��  	���A��*SYST�EM*��V9.3�0162 9/�2/2021 �A  �����AAVM_WR�K_T  �� $EXPOS�URE  $�CAMCLBDA�T@ $PS_�TRGVT��$nX aHZgWDISfWgPg�RgLENS_C_ENT_X�Yg�yORf   �$CMP_GC_��UTNUMAP�RE_MAST_�C� 	�GR�V_M{$NE�W��	STAT�_RUNARES�_ER�VTCP�6� aTC32:dXSM�&&��#END!OR7GBK!SM���3!UPD��A�BS; � P/ �  $PAR�A�  K\~�IO_CNV�w l� RAC��LO�MOD_T�YP@FIR�H�AL�>#IN_O�U�FAC� gINTERCEPf�BI�IZ@PO��ALRM_RE�CO"  � A�LM�"ENB���&ON�!� MDG�/ 0 $DEBUG1A�"d
�$3AO� ."��!�_IF� � 
$ENABL@QC#� P dC#U5K�!MA�B �"��
� OG�f 0COURR_D1P $Q3GLIN@S1I4$C$�AUSOd�APPINFOEQ/� �L A �?1�5/ H ��79EQUIP� 2�0NAM�� ��2_OVR��$VERSI�� ��0COUP�LE,   $��!PPV1CES00�!H �   A> ��1	 � $�SOFT�T_I�DBTOTAL_�EQ� Q1]@NO�`BU SPI_IN�DE]uEXBSC_REEN_�4B7SIG�0O%K�W@PK_FI0	$THKY�GoPANEhD � �DUMMY1dH�D�!U4 Q4ARG1�R�
 � $TIT1d ��� �7Td7T� 7TP7T5�5V65V75V85V95W05W>W�A7URWQT7UfW1pW1zW1�W�1�W2�R!SBN�_CF�!�0�$!J� ; 
2�1_�CMNT�$F�LAGS]�CH�E"$Nb_OP�T�2� � ELLS�ETUP  �`�0HO�0 PR�Z1%{cMACRO��bREPR�hD0D�+t@��b{�eHM� MN�B
1� U�TOB U��0 9DEV�IC4STI�0� � P@13��`BQdf"�VAL�#ISP_�UNI�#p_DOxv7IyFR_F�@�K%D13�;A�c�C�_WA?t�a�zOF�F_@N�DEL��xLF0q�A�qrc?q�p�C?�`ıA�E�C#�s�ATB<�t��MO� �sOE � [M�s���2�REV�B3ILF��1XI� %��R  � O�D}`j�$NO`M�+��0b�x�/�"u�� �����4AX�@Dd p{ E RD_Eb�~�$FSSB�&~W`KBD_SE2u�AG� G�2 "_��B�� V�t:5`�ׁQC ��a_E�Du � � �C2��`S�p�4%y$l �t$OP�@rQB�qy�_OK���0, P_C� y��dxh�U �`LACI�!��a���� FqCOsMM� �0$D���ϑ�@�pX��OR4@BIGALLOW�G (KD2�2�@VAR5�d!�AB  �BL[@S � ,�KJqM�H`S�pZ@M�_O]z���C�Fd X�0GR�@��M�NFL�I���;@UIRE�84�"� SWIT�=$/0_No`S�"C�F_�G� �>0WARNMxp�d��%`LI�V`NS]T� COR-r�FLTR�TRA�T T�`� $A�CCqS�� X�r�$ORI�.&ӧR�T�`_SFg�C�HGV0I�p�T���PA�I��T��� ��K�� �� �#@a���HSDR�B��2�BJ; ��C��3�4�5��6�7�8�9��2
���x@�2� @� TRQ��$�%f��ր����_Uآ���4@COc <� ����Ȩ3�2^��LLECM�-�MULTIV4�"$��A
2FS�ILD�D�
1��z@T_1b � 4� STY 2�b4�=@�)24�p� DԼ� |9 $��.p��6�I`�L* \�TO��E��EXT���ї��B�ю�22f�E��@��1b.'�B s�G�Q� �" Q�/%�a��X�%�?s��E�U� Sҟ�;A�Ɨ�qM�� � C��O�! L�0a��� X׻pAβ$JO�BB�����TRIGO�" dӀ���� �X�-'x���G�ҧ3AqC�`��b# tӀ�F� �CNG�AiBA� ϑ��!���/1��@À�0����R0P/pX����$
�|���BqF]�
2J]�_)RN��C`J`�e*�J?�D/5C�	��ӧ��@{ A�P�O�3л!% \�0RO0�6� �IT�s� NOM_8pn#�c� ���TU�@P�� � ��&+P���� ӨP�	ݭ��R�Ax@n �3�A���
g$TF3%#D3
�T��wpU�13�}�%�mHrzT1�E ���ޣ�#ݤ�%ߢ�QlYNT�"� DoBGDE�!'D�]�PU���@t����"���AX��"�uTAI2sBUFۆ��?!��1( ��P&V`P�I84'mP�'M��(M�)B �&F�'S�IMQS�@ZKEE3PAT�zЙp8"�"<!_MC��1)S�0��`JB�����aDECg:� g5�������* �U�CH�NS_EMPͲ#$G��7�_��c�;�1_FP)�TC�6S���5�`%��4�} ��V����W���JR����SEGF�RAq�Oaa #PT�_LIN�KCPVAFbag��`  C$+�� �ckBZ�PBzr�5,` +�ԦE� �A�0��Ad0o`Ar�D8���Id1SIZh���	T�FT�C�Z1Y�ARSm��CP@'�I c\1@cX�0<@L�����0�VCRCߥ�sCC���U1@�X�1��2��Mpq�U�1`�X�Q"�UDݤأiCk�p���
DK`݀f��RhE�VRf �Fha_	EF�0N�f�Pd1�&h���5�jC}�+�V'SCA[��A�f����4-)��p��SaFV�P#t1B L(�14��.�	�ׇ�MARG���a�F�@@���1DcQ���0LEW�-��R�P<���o�l:"RɄ/�������ȯ�� 5ڡR�� HANC��$LG5��a��Ӑ��ـF�B�Ae����0R�r��3@����@�@ ;�RA��@�AZ�0��N`:�O��FCT���p��F��R�0P0b ADI�O�a���a����&�ӄ5�5����Sp[�g���BMPUD�(PY�1��AES�CPjc�W��N  S~h�XYZWPR�cr����	���p}I��0  �P�I8���41��n@_�C�$ϑW�3U0M�MENU�2)�T#IT]q<�b�%ECAp:"�}���3 P�/EGED9�E����wPDT7�REMJ�<�AUTH_KEGY  �\`��  z~�Oa����!OERRLd��4�,&Q��OR�B$����z����UN_O7�>�P$SYS��4(������!qV�V@~pDBPXWO�Pz�5��$SKo��"��DBT�pT�RL�6 �C AqC����[�INDU �DJ�p�_�`�!X?���K�PL�A_2SWA��h�E��D!�u�!%RhM�UM�MY9����1� MMDB���7���!PR�Q1�O��9���8 г$�r�$ Q��LBֹ9����P�:	�^z�PC�;(�~z�PENEC0�TNr<G�z���C�OR"�=H �mO�@8$L��9$ֳ�"{���R@���VA��_D�� R3OS �"SK���Zr"��� =�ՠ��P�A��JVBETURYN���SMR(�U v#�CR��EWMDB=0GNALV �"�$LA� Y�*:{$P,p;$P��"�<m�!�PC���PDO^@,s�¯��R>��GO_AW����MO��pB��C{SSҐSTCY���>��R��0���IDT�R�2��2�N�СO@�J��v`I�� �?-�$L�RBl�Bt�PI�POj�I_BY,�r��T�VR=�HNDG��@ H�`�1_�@cS��DSBLI�����X0}�<�LS��A��0� ��FB��FE��~�7��=�5��=BK $DO�1�C"�MC�0o��4��7�RHɀW��K4ELE�Lr���ѯSLAVNrCxBI�NS ���#��=ᥕD�@,e��p񐳃
�{� 
��u��[!�٢BI���@�W��KNTV�#VE�$��SKIlA�C$;3�2UB�1J�f�1A�
DSAF7�5��_SVl�EXCL�U+���rONL��0 YW��Ȁ��H�I_V��RPPLYm�RysH� .�_M�O�VRF�Y_G�,M�s$CIOv0Ȁ{�P1UBd��Oh�1LS���N���4!��:@�P�$�ԄY�OCNE N�����,��GCHD���_����3ِAF��CP�c$TF1�A_V�AL�2[����� 3Em� �TA&��0N�p ��v�CLt	FxB�pT	��A<�P$�$��SG�` G� � 
$CUR 6�Sѿ���!7�?����(��&ANNUN�A��3�� ���� `�&�6931�P;:W6:��EF��IA�H @b�`F2���POTV� _㧴�������s0-M��NIݲI���2�G�0A�4DAY��LOAD^䜴�2z��5���EF(p+XI�Jm�%QP��O#@:�8�_RTRQsAK D�a��M@�yRYCE��bC#E �2J̐�wHA_����Afp=AqL 0�P1�AAyT�B,s�vD�UV��u��CAB2qM�2�`NS�A�PIDLE_PW�sh�EW��pV^�V_�@|@���DIAG��?N� 1$b ��ՓT*r�SrT� SZ�b�BRd��1�DVEр��SW�Q��
`��@D�HE@KVpHAO�H^E�APP�P�CI	R��BB`R�Ci� XҶAQ0�Rx��XP����U^��E@M̐M@���QURQDW�UMS�x�MeA�p�UxR�DLIFE�`Y3w`���bN�aTR�e31�cTR�a��32CC���Nr7�Y]pE�FLA*�f40OV��fHE�!>�BSUPPO&�M���bG�_ t�%�a_�X9�#t��.wZ+zW�+zC�.wу31��l�X�Z`�ͱ�AY2�xC"��T���RUN�0PU*31Jށ �V_���Ax}����O `d�CACH�#.��sS�IZ�f�`
^ғ�SoUFFI*p  }`�᜴B��6���!9Mq��tP 8?0^�oIMAG�TM����3l�8�g���D��2OOCVIE�PB�Qʒ⺰L|� 9?� �	 @D��tRU@6��ST� !Ԃ��܄��܄�0܄@܀EMAIL�0i�Y!<�^3!FAUL�2Sʒ,��-�AX��UԐ���$�A�T< �$G�n�S�@�@IT��BUF�9�(C����`Bs�b��C8��H��U�SAV����iP�rўPٗ��76PŔn����T��a_s���^!�OT����-#Pk��>��"A�#AX��t0vXs�S��_G�c
�YN�_�QC�U <�@D�i�M����RM�Bj�`T�F�$�6 DIY!�E5�I�$� B�V��"G���1�&�#��ˡ�q8��0F��� W (o�SV�У�����9�8�B�X����;�"�C_����K��k��"�f���Rd�e�,��D�SP|�I�PC��I�M˓��ɱ:%�b U`���`��[�IP}0I��Q�p��TH�p1�d��(@T����HS֣���BSC��p�@V� S�Q�j�Yğ�8DNV�G��YĤp��s�	F�Q��d��Ơh� ��SC3R_�[�MER|'�FBCMP'vH�ET�� YZ�FUpDUg���P�{r�CD��#�5�0�O �EOC0ɃZUC��!Q��RQ� Q�^!MAS,!/�N 2К4���?�� A|1[� �"�@�R��$ZO�L"���U4R���Pn��CNG����<����GROU��'B2XS�pGMN��L� ��L���L�P�`�����HR'�#����CYC�d����Ӥ�l���DE%_D�B�RO���$��T��0 ���410��3/���v �8���_�,�~q��A	L�p|1\��G��!��H�% B�Q����ERr7 T}Pʂ] ,��_�G�La�1\ �
MA�� �|1^�Ѐ$���5��EP�!��C� ������H���_H *LM/�# O ��U0 �zX!x��x�1xAxD�x7
u	8u	9u
�`w�
U1�
1�
1�
1�
U1�
1�
1�
1�
�2�
2��
2�
2��
2�
2�
2�
2��
2�
3�
3�
3T��
3�
3�
3�
U3�
3�
3�
4�&�XTDQ|1`��,�����֢��ŭ��'���  �FDR3T7aTS�VE�@=���b1QbRE��F���BOVM|�'5A�09TROV09DTlɐP:MX_<IN098�`O:0QINDn0pB!
�8נ����Gs��S�Y0��eyQD]FY0R�IV���ҷBGEA-R|�IOpUK 2�DNƠHwAnh3Ј���>�BZ_MCM~p�a,� �`UR��b�� ���? �`��?�l@�Q?lAE@�@tA������"c��j8`P��@PRI.����B�!UP2_� d ���TD�PP}�T@��A�G�E܍���BAC��e QTҀ����)�%�t\���nAIFI����pMa �P,UPT��R��FLUIǄ�f ��᪇I�UR a��b"�ޡQ�v�C�EMP����$�RS.\P?x�PJ����0�VRT� ��x$�SHO�QLob4�A�SS4�;��e��$BG_�
a+#
a�
ax�
a�FORC1�ط@gQ��g'�FUWA1ˢZc2�fR�p�L�h |�0NAV�����P�R�0S����$VISIl�0��SCK�SE�@��P8�gV�O��a$��0K��$���I@ΰ�FM�R2�%i   23г�1�v7O@O0OG6�0D5 2_�!��>LIMIT_</Q�C_LM�6�?>�=DGCLF�3�1�DY�xLD�A�45��6�?�4�!M� Ƀj���sy T�F9S�C�k P� O�|���$EX_O��f�O�1g�����O�3���5���Gm��%l� ��0��SW��OyN�V3EBUGdL݁%5GR@୰U���BK'�O1J C@POWp�����ǅ�M��OV��S�M��E͒�A�0��_?E m m`��/TERMX�na���'ORI�]�oa�D`KSMc�O�B]�pa����Р�qa�� �U�P<� r� -�1��m�Po���n�`G��pELTaO}Q��Ѡ��FIp��СW@Ӂ����o$wUFRR$��0�J�ՎpOTW���qT2�0i�NST���PAT(�}�PTHJf��E��(����ART�p���p�w�"�REL��'�S�HFT������_��PR��Ӟ� ��$���q�qp�P�㢡R��I䠫tU ПPAYLO����DYN_iP�@�R��za%�ERV� P��R  ��"e�����!HP���+!HPRC�AAS?YMFLTR�#WJ(��!�0E�C��۹�R�U����`������ɥP��j���/�kOR��Ms��G��$sUb�-���D���L�H��C�t ԰k�LU�`3�OC�|���$OP�d�����S1�P��RE��R,���_�h��e�PR�����|ˡ&Te$PWR�0]�c��R_�è��`c�"�UD�B����5�w u�@$H%U�!��ADDR��H�J�G���ѠљѴ�R��b	Qv H� SSC�b#��+#�՛��ƨSEC��c��HS�CD_MNmRw��`��2���r�HOL}��"���%�&���CROy`��QND�_CG����^�T�GOROUP����_y@�b���1t
2�� �� ��%1�� �� ��� 
2A�`�2��SAVED��%����b�#�P�@��_D� H��R�P���bG_HTTP_��H	Qwy ( OBJ�`l��&T$��LEv����z�
Pz � (�'�P� _�1T=���qS��A�xXKRLH�?HITCOU1 ��QL�a�����R�V�S���JW��SS�0�$J�QUERY_FL�An�߰_WEBS;OC�b�HW���	Q{��e�INCPU���aO���_`�˃� �ԣ�ԣG" ��IOLNR| �8� RP�`$S�Lg�$INPU�T_&q$��Pn�c T� SL&�
	Q}� �*&³��²~�IOY�F_�AS5�~P$L�P��#Q��aZ�,�`�P��P�R�HY�'p����]UOP2� `n���~2�~0���PA���@!�"&�`M���nQ� ln�8�TA4h���A��TI%+Ű�PWpi%ϠPSh&BUWpIDG����%����%@�7"�"w��D!I*|$]$� N�(�Wp�%�IRCA_�CN�  � �ھ�%CY��EA �1�a#<~0A�;7�S�l����#5�DAY_<� �(NTVA}U� �7���#7SCA�b�7CL�1�!�Q��"�`nQ��/�$���%�5N_��CNR� �"m1@ �!L`��/A���� �!]�s8La C2��@6#&QnQ�R8fF��f LABw��A\Wp�GUNIPQxC��ITY�8!���R!R3���҅PR_wURL�`�$A3�EN����a��n�T�]�T_U�TABK#Y_2`:�~�J� nQ� X� 'Rߵ�Q� R�HP�pAӄ$RQJ�R^QFLq��P/��
qS�s
�UJR.tň ���Fy�.���PC��RD�3$JY7��bJ8�Y7��Hr2�R�W7�F�P8�Y��QAPHI�pQ��SgDc�J7J8��0`L_KE�@ � �K� LM��! � <�0X�Ra� 3WATCH_VA�am��A��_FIELD��yA�LLb2�� �pm�VZ���aCT�@�f[���� LG�C��� $9LG_SIZ�����e0��fe�fFDxI�hx)�v �hZ�wx�`���c|v 0�|ve|v%p|vZ�|v�˱ǅ�_a�_CM [��qx��z�qF��w��t�`�(�a � q�p�e�%p&�I�0�)��Z�2��$��`RSo`��  >�ZIPDUQ#�1SLN�Qw� DE�qE+;`���A�a�Á��L̃DAU�EAi�� ������GH��bAqBO�O���� C�=pITN2��ЄsRE> I�SCR����D���MARGIK�}�	|��ħ�qS��pWp��qׄ|JGMݗ�MNCHn�qFN�Bb��K� P�UF��/��FWD�H]LI�STP�V���@�9��RS��HG�.�yCY�_���|I�ݩU`�&���z��Ǖ�`��G����P�O�d�t�_��r��O�C�B�EXxTUI�IUpC0Uq�� ��Γ����A$���2�e���e�NY�n�AcNAq���2AI�P8_��3:UDCSp0�Ө����O�O*�S�SH�5�SAȜ�IGNp�0 s��`>A!�7DEV��LL<Q� Hq�2@ ��`�!T�$w�H�4�Q_�-A����`�0� ��G�$8�1�2��3�HaM��@ �# ������H� ��%I�L8�G��Q|�+ST�R��Y:�ѿ �$E��C �ۼP_����u�M��a� L� ��p�� ���0��_i�0��a���e�_ �b@�� n�3f�^��M�C��� ���C�LDP�:UTRQ�LI�A<V���FL R�I���1D�a���v LD����OR�GBQ�����xRESERV������q�S� � �	�帥���mpPT���xR	��m�u�RCLMC���%����� u�c@M��`�@��Y`$DEBUG�MAS�i0ZC�rUR��T���%E�PT�����FRQ�� �� �iHRS_KRU(�1DA?0��FREQ�p;�y$���gOVER~ � s�`J֢VP�EFI� %�2D����9@�� \2PS��T$UP�/B?�J�1PS�]P	�^C���X"���U|� ��?( 	�Q�MISC�U� d���P�RQ[R	/`TB���  G��T�AX:RG`WpEXGCES�B/�*M  
�A�� ;:T��*;SCQ� ��@-@K_]@ER0�n�/��MK�D���R쐐��B_�`FLI�C�BS�QUIR-EƣMO:,OJ+��� ML*�M�E� �X�A�� �b(#��F8�NDԁ{0  ���ȴ��h�#D�sЄIN�AUTv�ЄRSM�P�(m�N�Ҕqܣ�!���!PSTL�A�� 4�0LOCS�R�I�@S�EXH6ANqG���ODA#��7�B�P�MF�b,u�y�)⃰3帳5����SUP<� � �FXUPIGG>E� � �)� �q)�Ц)��@��� �9��H��F�:������TI�`	к�p�MEP�� t{0M	DxA�B)�F��D���GH\0�Q�DDIA�Q�CXPW���D��m�*�ED�)�O�Smpn  � �CUp�V�@e���O��_��Q� �}�[Ӆ3L���0pBXPB^h��d�IPPAXKEҢx`�-$B�5V'��ND2��tc�Q2_{TX2�XTRA�4�R���� LO �  1���TC�V���	R�V�S�RR2>.� 0�Q��Ar� d$CA�LIM�uG�0g2�Jh�� �RsIN�4c<$R>`�SW0��c��ABC�8D_J�PA!P��A_J3�f
�b1#SP; �@PP�d�m�3�mQ��P�eJP��u4�lqO��IebCSKP��:t�p$�:tJ�Q:|kupQukuawQ0_AZq�q�qEL��r��O�CMP_3�ȀR1T�s�U1�p�UFs�1��x���zZ�t�SMG��i@��JG�P�SCL�L5SPH_M�]�>��@P=;`RTER`4cIܰ1`_�_�x�aA����{�DI�qn)�23U<rDF�0���LW��VELƒ�IN>⨰ŀ_BL��̈́fbJ�҇<��MECH�®�OTSA_a�0!1#IN^�S  �	R/�П�Q-���_ ��<�W���� T���a����0DH��P"a���$V=`�#7����$�iDd��$���R�C  ��H �$BEL��p3[�_ACCE�Ӂ �����IR�C_|�7�NT<�}�$PS���L�0P0C���/�$� �1�%��Q�z��z�3I�@�_�Β��p��d� �_MGCcDDΡ|�DFWu��j@
����ߨDE��PPABNQ�RO?�EE���8����aq�����'�$U�SE_<`سP�C�TR״Y*���p� &�YN-A�p��*p��A��M Q6ȠO8��l�ŴINC�DY1���T�faUENCl�LPA�A��R>�IN��II�.�k@�'�NT���NT2c3_��D\�LO��Dr�{ I� �|Ʀ�@	�	�0���CG�C�MOSIӡ"!P���cPERCH#  
�ya� ��_1 ��2A¼�2A�w�r��H����(sAI�;�Lx� (s�'wD��0�z֕�gTRK_��AY�S 5����I��ծ�Z0�v8���� MOM�BT@�	�P��0g�Ә|�]�`DUe`��S�_BCKLSH_CI�<�  ��z ����[��e꯱cuCLA�LM@��Ѐ���C�HK=p\@�TGLRTY6@�S.�]E��iA9_�3��_UM�����C��ܡ2��G LMT�`_L̐�s��A&�E �A�3��6�<��6��`��D҂��PC����H�0h ҥ��C�MC�Uܠ�CN_bKbN�S��sSF��V��[A$�[���I��%��CAT��SH �3Kb����%�%��U0J��Y�pϠPA���_P����_>p2���`��=q�����JG�0�����OG��g�TORQUt��e������+"��h��8_W ���qϑW��VƓ�VI^IlIƓF�r0Ir�!qؠVC"�0���1�Р8��q�JRK�",
&PDB0�M:SP�M� _DL��U�GRV]V$��V$Ɠ7!�H_�S5#}��*CO1S�+�p�(LN �+ ��$���)��)��*��,�2%Z� ��7!M�Y�!08�"�Q�+Q9T�HET0��NK2a3Ɠ{2��� CB�6kCB��C@`ASQA��2��1���1�6SB8���2�5GTSCqP�C�a��w��wJ�#$DU��^�,Bab(ԅ;G�Q�_��n+NE@ti�K���y����o1As5�E�G�%�(�!LPH�%zBT�zBS��C�%�C�%zB��&SZ6�@V�HV��H���LV�JV�KV� [V[V[V*[V8YH�H�F�R�MZ�X��KH [H[H[H�*[H8YO�LO�HOTii�NO�JO�KO [UO[O[O*[O6�FzB�1�i�%t�GS�PBALANCE�_@1,sLE�0H_s5SP4��&Tr�&Tr>�&PFULCXxr�gwr�%A�1��qU�TO_����T1T2�y �2N���L� �t%��сp_@P������Tk�O���GIN�SEG���REV8���=�DIF��f��1�K���1���O!BA���`#�2"L����?$LCHWARL*���AB������@0����X��P�e�ֆ�G���p� 
pׂ5��&�ROB���CRC����	���C��_�T �� x $WEgIGH����$�CdR�� I��z�IFl�N�LAG����S���0���BIL��OD��С�i�ST�i�P0���j� ސD 9�B���F�

������ � 2���n�DEB�Uz�Lr���+@M'MY99�/�N��΅�$Dr���$��� b1 ��DO_0�AA�� <U�Ԗ�p�A���@IB����N@�w�_��ꦰ���O�� �/� %	�T-�5���TB���<�TICYK{���T1D�%̣�3�ՠN���pk���R�R঱��祟��K�P�ROMP��E�B $IR����8.�N�m�MAI< ��4��G�_��E�N�t�Ѹ�RK CODٓsFU��w�ID_�����.�(�4pG_SU;FF� ���N��DO�%�����GR����Ǵ� Ӵ��޵���AǴK��㐮U�Hu�_FIvؑ9=�ORD��3 H��36i�>�|��D�$ZDT�������N��4 *M�L_NA��ՠ��>�DEF_I�ȗ� ���󥫒榵��������ISc@ c�r@�&����,
�4��|�D�p5�\��ٓDO6pb�LOCKE�������(�ǲ��UMƵ��Ǵ ��Ǵ��Ǵ4�Ӳ��ҵ ��Ӵ��Ӳ��(�(�޳ ���޵��޵��޳/�m�ø��Ps�Ԫ�"�Dx@<�W�ا������TE��O��(� �LOMB_t����0i�VIS� WITYi�A�O��A_FRI�s�t�#SI"��daRҠ-��ݠ-�3�i�W	�W��G � _x��EASq����r n�TM�.�4+�5+�6r��ORMULA_I����THRq� ��G�ǲF�y0�8��COEFF_O ���/���0Geq�Sz�+�CA�p0�B�a$��p���GRc@� � � $h���rl�X��TM�����տ����u�ER�?�T�Ԇ�7��  ��rLL�f�S�A_�SVa�����7���$07�� �SwETU"�MEA=�����j���>�B�� g� { 
� �����B�vэ��Hՠvђ�s�cZ���o�=�n��tQ@v�a�RECQ�z�H�MSK_7pޏ� PU�1_USER�q�2$��8 4 �qVEL� ���C"7%��Ip��p��MT��CFG!�O  נS�Oł�NORE@���"��OPWOR}@ ��,8�SYSB9U�P�SOP�! J�T�*U�+N�P��a"�%PA ��#��V�OPܰUw��!�s�֒�0IMAGd��p0Z�IM� �25INx�223RGOVRD\P�# 1P013�r@]�b�5�ƂL��BTqB�P�MC_Ex��!�N"�`M�2��1�4��^1SLrp � � $OVSL�S��DEXR����5W@��>_^0G�_0�C�C*G%H�JCC�����5YA'G_0_Z+ER�!�3Mx�Ɓ�G�4Ł �2P!�O @ uC��O��RI�A�
�F]��I��A�A��P�E]A �� HU���ATU�S�"�C_TI1DXVB� VQ�L�p��Cx� � DY� 0�CQ�P#�QC�3 ��1XEP�kRR�JT�C��@V�PUP�>��PX1�=V
A�
�3�7FR�PG�o%�� $SUB�Q��
�Q�CJMP�WAIT�PCeL�OWłF���FRC�VFU�ؠł aRE�Q`F&���C\@RL�łؠngIGNR_{PL�CDBTB��P �ƁBWu�dd� U��ceIG�!��q�ȀTNLNbf�bR-T�3NO_�N��3�PEED�P�3HA�DOW��ă� ER�VE�3t
B�Q��S}P�p � LU�`݀��1p'�>tUNg���[=p�QR�PdCLY�m��Q���9Pb !� 0�@�"�2�O�LE�Qn�P�A�Є����f!PI�P�b!� h ?$ARSIZz�D��3����@O�9b��A�T���c��r(�EM2τ�tcsUX� pB��1PL��p$� $z!��SWI��ł;��WO���A��?�L�LB!�� �$BA�DlӴB�AM�@$�C���AF��J5-p�q��6��>h�_KNOW�sςb0U�AD��i <p�D �PAYLOA����_Q��!*�Z�L
�A����LCL_�  !�JS���U!`�s2
n�Fx�C� N��Q�
�IN�R� N�ߑrP2l�B��� _J�bؑ�_JX�6!�PTAND˒���X�l� ���PLu�AL_ S�L�<pA�B�1���C�D�E��sJ3��� T�p�PDCK�0ҴC�Oc>�PH/�u�BaED�/�A��^|�a�0 � ��`��D_1�2A�DcARrQ�ߥ�lPRTIA4�5:�6�MOM��)��I�6�I�C�l B4`A�D)�m�6�m�C�PUB@RN���6���C���q���ܑ~�� � �pM��`Y �'r@�$�� e$PI�4�aΣ'!�P�SA6��I�I,�I:�ڴR�k��Qk��Q$ROk��C��E�cHIG[��c5e.t ��.t5ek```�������ka��ka5eSAMP zP�q!ٴ�'�5e����  U�� t�7" d��Pn�.p�}��7"�R��"�lՅ���l�IN�܅�
Ӽ��۳�5b���������GAM�M��SQ�r�BET���FI�sA���T"
&]IBL�bIƀ�sO$HI���AP7"��E���������LW��������栮�^���`!�C�eC�HKl0�@�d�I_	Ќ�U!��̩�р��h�I�g�g�� ��$Q� 1��k�IRCH_�D%#��PVd�LE@Q!'!�A��������`�MSWFLedɱS;CR�X100#2 d�e�J��� )�}�x]	.plPI3A�METHOpC��eV�AX�CwPX�`����bERI�&�3�R�RQp�	����FH5$'�k�z���L��'�)OOP�k��?z��APP�cF�0�pCdO&��RT��O
�.p���pR۴�@1��۴S@�:��RA��pMG�a�r�S�V}��PS CU9R/!GRO�`�2S_SA���4!%�SNO��C�A�R��!  q�̯"�4�@Ȏ*~+f���nŻ(�DO-qA n��`d�_
�ծȸq�� �q��75�#W�n��@:?�M�� ��0��YL�̑���S ˒"�Qq77͑(��}3̑_��CraiQ'M_WP �2/��3+My`�;s��7��Bd8t�7�R�M�!�B� � $�h1`B�QW1@�$�L�AD�1@��/B��@/B��/BC��`��N�pPs�R����XypO�����Z�E�?`�� ��M��f&c/u/��/�/�/ ����uL:��_�R� |b��H . I�{V6�{VC�. "�`�W�V<�a�k� 鳜_R�� װ]VP��q�PMON_Q}U+� � 8�p�QCOU���QT�H�`HOj2&`HY�S�ES��&`UE�`"�pO�t�  �N�P@��B!RUNW_TO�3r�O��N�� P�oeC�1�>� INDE�R�OGRA�06�~02>�0NE_NO�doe�ITⱽ`S`INFO�Q� N��j�a�|2�O1OI�b� =(k�SLEQ��q0��p�f-@OSA��t�� 4�pENA�B]Bm`PTION<�s�PERVEs�jw����BsGCFKqԋ @`J�0��wb�w�R�xk}wYR�ΰEDIT�Q� I�>@�@Ḵ�����E��NU�w�xAUyT=!�uCOPY̱P�����I M��N ��$�9�PRUT� �'�N�pOUC���$Gtb�YRRGA�DJ�Q� hb�X_�0I��@���@��W��P�� ���Û�z��N��_CYC]B��RGNSGuל_0) LGOF��NYQ_FREQ��qW	���<�SIZZtG�LA�3���D�	����CRE~�G�I�F,��cNA/�%�z�_G�STAT�UbP�egMAIL�-�q�ő��!dLAS�Tőp��ELEM�Kq� �H UxFEASIXq2Z�S F ��*!%����}�I �`{�3���)a�P��Z��ABAa��E�`��V�r�BAS��s�}�ⲱU����6 $,����RMϰRT��р��£�C�������� ������jP	~1� 2� �� �D�������@���1��B�
���DOU��c��^�P���ڞrGRID�aAcB7ARS��TYYsO1r��O�P�Q� `aE_��!׀��}�O�@>Ht� � �0�P�POR�c泗�S�RV��)���DI? T_t� �2ā�<�T��<�4:�5:�6:�%7:�8��QFN�Kq��^`$VALU���%���FGu�� !TuJA�aг1��(� AN#��𬑈@��TOTAcL_ɔX�"�PW)��I��7�REGEN5�J��SX���c)��Q���`TR����5�_!S ��J��V���t�҂rs�E̓� +a��ob���V_H��DqAS����S_YE!��BM�S$@ARP2�� w�IG_S!E"c����ܕ_s`��;C_��$CMYRE�c�DET +�q�I�I�Zb�<㶲��ENoHANCa�jP�
Tw��P���IN�T���0Fic�AM�ASK���OVR��`� (P���q��OCVCf����È��Pr�6�s۱��PSL�G4���� \ @"�FB�ʐS�2ݔu�UEeg����Ӥ�F�U P0o�T�E�@��� (�rѮJN�="]�IL_M\� V`�� �PCTQ`��a��C�Vj�2V:CHP_ �6 RMi	V1h
VU1v2�2v3�3v4�4v
!C�� (��1�"INVIB@B/�!�6222>323
>424>�PQ^R M S�`�vPL��TOR`�%IN��#m�."[0��d�0MC_F,/`D 0L!!���MN I��""^�� lPRu��0KE�EP_HNADD"!!]$w�g)C�A��A}$��"��~#Oa�\$*�!0~#��~#REM�"}$ɑ಺%��!�(U��e}$HP�WD  ]#S�BM��װCOLL�ABD����р���`IT��@5�NO�QFCALTC�D�ON�l�"�D� �,��FLZ@��$�SYN �<M�PC�O����UP_DL�Y�Q�^bDELAh�0ʑ��Y�PADQ}��QSKIP3E'� ���q`O@��C�0P_q`�bG�` �BՀG�q+I�q+IS� *J`�*Jm�*Jz�*J���*J��*J9U��J2�R��@�PsX��T 6��A�a��A��Y"�A8�aY!�PRDC��2�� ��pR�s�R�o��)b��RGEp�pC��g�FLGa�(0��SWgy�SP9C�c��UM_�@��_2TH2Na��P~�@ 1� �@�ED��Gr � �D�`��eY{�2_P�C��RS��֡=�L/10_C[���U�� ꣀ}�6��  ?U�C#aT�q&:��Q�Vc�`���H�{�H��V��P� }P�PDESIG�R.6�VL1�Y1�Vscv�g10� _DS�Cr1��/�11q� lN �!�� UsA3�AT� ��l�?�rIND����q/��q<�r�HOME<r
�
�d2�b��o((:L�g3�b�o�p���� ��d4�b����"�4��F� �d5�b��i�{�������Ï�g6�b����
��.�@�
�g7�b�c�u�����(����^w8�b���� ��(�:�^uS!0�a�  ��c_��aP�c� E�� aT�P���IO����I��D�O]0_O�P�6��� �$�ASSaP��i�c�`P`P X����SI* a��n�1r�$AA�VM_WRK 2� c� �0  �5�j���ĸ��� �	�`���`Pd�!��I�0�N���m̀y�	�ϴ����Ē�B�S�pQ 1���? <��� %�7�I�[�m�ߑߣ� �����������!�3� E�W�i�{������ ��������/�A�S� e�w������������� ��+=Oas ��������'��C�0AXL�MP�*���  md<INE�S�;PRE�PEh��w_UP-b���c���IOCNV_ԋPH�SP�US؈����IO�0V �1��P $���`4�-��/d�?�* J?/Q/c/u/�/�/�/ �/�/�/�/??)?;? M?_?q?�?�?�?�?�? �?�?OO%O7OIO[O mOO�O�O�O�O�O�O �O_!_3_E_W_i_{_ �_�_�_�_�_�_�_o o/oAoSoeowo�o�o �o�o�o�o�o+ =Oas���� �����'�9�K� ]�o���������ɏۏ ����#�5�G�Y�k� }�������şן��� ��1�C�U�g�y��� ������ӯ���	�� -�?�Q�c�u������� ��Ͽ����)�;� M�_�qσϕϧϹ����������%�<LA�RMRECOV ��nw�LM_DG ' �*}�_IF +X*����������9�K�]�o��, 
 ���$�@0,��������$�� :�!�^������������5NGTOL � � 	 A�    <PPINFO �� ��EWi{n  ��}�lҚ �����.R<b������� ���/ /2/D/V/�h/z/�/��PPLI�CATION ?}���u�Handl�ingTool ��% 
V9.3�0P/20 �'?
88340�#�*7991029>�231�%�*�/�"�7DF3� �,�#N�one�+FR=L�/ 22=�&_ACTIVE2�s  �#��  �3�UTOMOD�0�����5CHGAP�ON�0�>���0OUPLED 1��� 7@;OMO_O�;�CUREQ 1	���  TiIiL�iL	�O�E� �Dm�wiB��%ƯDH�E:B�JHTTHKY�OnҜO �O�O�O8_J_\_�_�_ �_�_�_�_�_�_�_o "o4oFoXo�o|o�o�o �o�o�o�o�o0 BT�x���� �����,�>�P� ��t���������Ώ�� ���(�:�L���p� ��������ʟܟ� � �$�6�H���l�~��� ����Ưد���� � 2�D���h�z������� ¿Կ���
��.�@� ��d�vψϦϬϾ��� ������*�<ߖ�`� r߄ߢߨߺ������� ��&�8��\�n��0����L{ETO���?��3DO_CLEA�NO�4>�NM  �� iO����������oNDSPDgRYRE��5HI�0h�@y�@Rdv� �������8MAX� %����AG6X%�512B51�2PLUGG%@&�2C��5PRC��Bf�"j�/!�O� ^SEGF�0K� ��f�x�@/R/d/v/8�/��LAP0. �C�/�/ ??$?6?H?�Z?l?~?�?�?�?�3T�OTALX��3U�SENU *K ��O�B{@RGDI_SPMMC�]�C!H@@*DO� =%&C_STRING 1
�;�
�M�0S��:
�A_ITE;M1�F  n�=�O �O�O�O�O__/_A_ S_e_w_�_�_�_�_�_��_�_oI/O SIGNAL�E�Tryout� Mode�EI�npG`Simul�ated�AOu�tYlOVER�R  = 100��BIn cyc�lMe�AProg� Aborcc�A~CdStatus�C�	Heartbe�at�GMH F�aul�g�cAler�io,>P�bt���  !�K!�O���� 1�C�U�g�y������� ��ӏ���	��-�?��WOR��Kw�� Q�����ß՟���� �/�A�S�e�w�����୯��ѯ���PO �K�a����>�P�b� t���������ο�� ��(�:�L�^�pς����DEV���2� ������
��.�@�R� d�v߈ߚ߬߾����������*�<�PALT�}cᏟ=��� ����������	��-� ?�Q�c�u�����������Q�GRI;�K {���/ASew� �������+=Oas���0R �}�����	/ /-/?/Q/c/u/�/�/ �/�/�/�/�/??�PREGg�P0�)? w?�?�?�?�?�?�?�? OO+O=OOOaOsO�O�O�O�Om�$AR�G_w�D ?	�����A��  	$�f	[X]W��g3Y�@SBN_CONFIG,`�KQa�PbjQKQCII�_SAVE  �dsQfS�@TCEL�LSETUP ��J%  OME�_IOml%M�OV_H�P�_�_R�EP�o�JUTO/BACK�Q�ImQ�FRA:\�=; 'o=6sP'�`�`=7ph� ��klP 2�1/11/23 �18:32:24=64X==�o�oal��<cu����=6�Q��� !�3�E��i�{����� ��ÏՏ`�����/� A�S�ޏw����������џ㟺�  \a_�?c_\ATBCK�CTL.TMP �G.DG GIF .T
/�A�S�e���V$sf�9cI�NIf��ecV9cMESSAG�P��sQ�PeSwQ��ODE_AD�P�VcU��ʢO���ӯ9cPAUS/� �!��K , �	�4P�E3�A�,		+�e�O���s� �������Ϳ����=�'�I�s���TSK  �po*o<`�UPDTʠ��d����XWZD_E�NB��_Z��STAp���A���AXISQP?UNT 2�EpQ�rP� 	 �GP �&�f�� ��P 1�. ��	=:nK�  
mPP�f��  5 � �fߟ߱�s��Go <>� J�� "Q� ?,� Q�����p����%�(�MET��2�ƏS PJ�D��B�D���D��
�E%^D��oEI����<a�<��r�=.1�<�l��<�;5<����.�SCRDCFG� 1�ERa ��UpR����� ��0�B�io=:���V �������������S� w�4FXj|�0��/�G?aGR2���X����NA�P�Ks	?d�_ED���1��� 
 ��%-�EDT-���[BG_LOG�ICK�
����P5@b>=:4R2P�V7����2��[/;/��P�@a�	/t/��c/��3p�//�/@/� U+��/@?�/�//?�/�4 x?�[V?�?��U+�?O S?e?�?�?�5DO�? �O�?�>mO�OO1O�OUO�6_�O]_�O�>�9_�_�O�O�_!_�7 �_L_)op_�>opo�_�__o�_�8�o�/�o~<�=�o<�o�o+�o�9t�o�?�=��Oa���CR�o����Mm g�ҏ�+���O�� ?NO_DEL���GE_UNUSE���IGALLO�W 1�	  � (*SYS�TEM*�	$SERV_GR!�܌��REG��$8��쌐NUM��ߓ�͝PMU8���LAYD��?PMPALt���CYC10�,�x��R�ULSU�0Ν.����Lh����BOXORI��C�UR_��͝PM�CNV���1�0B���T4DLI�������	*PRO�GRA��PG�_MI�D�V�AL($�c�M�V�B�����$FLUI_RESU2���ğ޿�#MR�������� 4�F�X�j�|ώϠϲ� ����������0�B� T�f�xߊߜ߮����� ������,�>�P�+��LAL_OUT �{���WD_ABORt�\�����ITR_RTN � �t�e���NO�NSTO�� ���CE_OPTI�O��g��ROIA_IY���$��h��FCFG ��
%�~M�_P}A��GP 1W�i�����������C�  �� � � � �� � � � �z � �  D��+DB B ���Y� � � �� �B ��D� �DB  � ��D3ʆ =B F� DYe��v?� �HE��ONFI����G�_PԠ1W� $���"4F�Xj|�KPAU�S��1�D�  B�~����� / &//J/\/B/�/f/�/��/�/�/�/�/?�M~��NFO 1��g� � �	��c?�pQ0B� ?�`  A �q�� B% �{ ��7�D��\D���A�16(�C��0�?�6�OQ��W��w-�OLL�ECT_Q�?6��f��7EN$����n�3NDECG����1234?567890oG�r঑g�mOF�s
 Hp��s)�O�O���O�O $_���O_h_3_E_W_ �_{_�_�_�_�_�_�_ @ooo/o�oSoeowo �o�o�o�o�o�o�`+IF��2K� M KMBIO  XIA���������wTR��2!�}(@��y
A&�� �"�}P�]� I_M�OR�r#��   2C4�مP1ى� ߏ��9�'�����q$��,�?�� ���@�K��?��P�2&O��������d�
ӟ8��7a�^��d�@j��5B�d� �sja���PDB��(��Otcpmidbg���ޯ� �:�E~šp�ʯ#��I �E~ȯg�2�5 F����63��mg����ĿF�f�A�=F�Spud1:fϏ�k�~��DEF '�(��s)z�c��buf.txt��講�.��_MC��)��sQd-�Ӹ�*ݤd��[�>�A��Cz��0�Ay0C7�B��wB�SwC�3�C3�C����l=D@�C�}�C����D�g�DM��EB�l=E����E�\E����F���F5ПF��-��1� Q ���b�,�|8��7�A)�@�N��Z� �d���px��L�ѥ�Cf q�Dր�$D�j?E�H��D��DA F���3E F�I3�l=FF��E���EA H�F�A G������ ? >�33 ���n��m��5Y��m�)�m��1��?�=?L��<#ס��q�|��O��RSMO?FST %��?^,6P_T1�s-�}�A ���MOD�E .����XY��1;��9��3�?���<��M>�̼��ES�T��+���R	B/��?c_�ՁA����D�0L��1pҒ C�@�B��Ck������0:dڡ� ��P1�	��*HIQC0R?g��1���D8�RT_~��PROG o��Z%��xE�pNU?SER  8E��dBIKEY_TBOL  ���J2��	
�� �!"#$%&'()*+,-./xG�:;<=>?@A�BC��GHIJK�LMNOPQRS�TUVWXYZ[�\]^_`abc�defghijk�lmnopqrs�tuvwxyz{�|}~��������������������������������������������������������������������������R!���͓���������������������������������耇����������������������qLLCK�Z���STA���/H_AUTO_DO5F9Y3IND0D�.b�1R��?6T2Y?��STO�@@?�0T{RLNLETE5G��:_SCREE�N ��k_csc �0U�0�MMENU 12�� <gf.O }O7OlOV�IOoO�O O�O�O�O�O_�O�O #_\_3_E_�_i_{_�_ �_�_�_o�_�_Foo /o|oSoeo�o�o�o�o �o�o�o0?x Oa������ �,���b�9�K��� o���������ɏ�� ��L�#�5�[���k�}� ʟ���� �ן��H� �1�~�U�g��������ï��ӯ�2�P��3R�E3�ɩVvq��EB;� BB�7B6KSW76�9L���0_MAN�UA���?�$DB;CO70RIG�7�)���_ERRLT	4�	��� �2�� ��NUMLI�Mz35�ZDB�PXWORK 15����Ϥ϶���|�� �DBTB_�1G 6�[ӯ�a���DB_AWA�Yó	GCP rZ=��.�_ALP��/.ҿ�Y�0�5Z ���_ݰ 17�� , 
�θ5�2s���,����_M60Ik�<��@��ONTIM6�7�Z�$�z��
���MOTNE�ND���RECO�RD 2=	� y�����G�O��������=�XECUTING
���	�� ��$�K���o������ ����-���Q���u� <N`���o� )��q&� \����;Q� I�m"/4/F/�� |/��//�/�/�/�/ i/?�/B?�/f?x?�? �??�?/?�?S?��� O(O:O�?^O�?WO�?��Il�O�O�OLO_ �O�O7_�O[_m__�O �_�_$_�_H_ b�o o(o�_Lo�_Eo�_�\�o�o�o7o��TO�LERENC;�B�Ȅ�I�L�ͻ�C�SS_CNSTC�Y 2>r��1��o���<J\n� �������� "�4�F�\�j�|���t�DEVICE 2?'{ �ޏ� ��)�;�M�_�q��������sHNDGDg @'{w�Cz��|��qLS 2Aȍ���)�;�M�_�q������rPARAM B��kҪ������SLAVE �Cȝ��_CFY�D�����dMC:�\pL%04d.'CSV��T�c<���6qbA i�CHq�ڑ��ߕ�|���ǧ�gࡲ�a޿̹�S�J#P��S�������RC_OUT �Eȍ�љ�_NOC�OD�F����S�GN G��z�#�M�11-�JAN-23 1�2:37l����23-NOV-2?1 18:4��� Sw�
������������M��Þ�j�������VERSIO�N ��V�4.2.14��E�FLOGIC 1�H'{ 	�h��������b�PROG_ENBo�Ж��WULS/� ϖb�_ACCLIM0�������W?RSTJNTO�y���b�MO��v��0�INIT I'z��� .�OPT�� ?	m�F�
 	R575��V��74��6��7��+50��1��2��h���\�}�TO  Љ���C�]�VT�DE�X�d'Ⳁ-[�P�ATH ��'�A�\RAC21-�CLUTCH-2�2.03.202�3\I����eHCP�_CLNTID y?@��� �o� ���bIAG_G�RP 2N� �qa 	 �E�  F?h Fx E?`RD��D 
qobl�p��Cfu�}yu�Y�dCu�q�B�i�	�mp3m6 �78901234�56�?�C � � A�ffA��=qA�i�х�A��HA�i�����A����"�@�i�pXi�HpA�ppl�BV�"���"��
�(�A�A�
=Aޙ���A��
A_�Q�A����i�@Rdi��xi��{A�J��Ʊi��_���A�-���Ϳ���/��EG�A@i�:��RA5� /)*-#�� � ���K/]/o/�/�/�Pz��AJ�!?9�p�A3\)A,/��A&Q07p@�/�/�/??�c�_]��AWQ0PU0UJC<�4U0-� %G�c?u?�? �?�?�7M_OqOOO�O �O1O{O�O�O�O�O%_ �O�O_m__]_�_�_ ?_�_q�D �4!�!�L1�0_=�
==��G�#a>�Ĝ�+e_7'ŬGe6�7�Se_@ʏ�\of�p�{e��@f\Ahi��`A�i�<i��<xn;�=R�=s���=x<�=�~Z�_;���e<'��g�� �?+���C�  <(��Uǲ 4kb���v���#u	�!��?g�_Y�]g� �k�t��o����/�A��Y?)7L�?S�Fg�$�/do�_�$`��G�_A�al�A��_L� x݃A�凯��C�0��@U�_�B|��ED  E��  Eh� D�������ܟ"�<��  �]�����	������Gᷤ���?f���?��6����6�7D�?��D���'���@ʟK�Ɵo�"���䑢	��:ǟ�j��@�e_��[���(���L�7� >�"=�"����ܼ��������U<����;ě����CT_CON?FIG O{��ßeg��!STBF_TTS�
����7���D�
��l�MAU��j�M_SW_CF˰P.�  OCVI�EW�Q^�j������������
� �Ҟ�3�E�W�i�{ߍ� ߱����������� /�A�S�e�w���*� ������������=� O�a�s�����&����� ����'��K] o���4�����#��RCW�R�U+�!��[��������SB�L_FAULT �SNs�!GPM�SK �)'��TDI�AG TϹj��3��aUD�1: 6789012345�"㲤a�/PI��/�/�/�/
? ?.?@?R?d?v?�?�? �?�?�?�?A�v&�	<r�
�/*Ou�TREC	P_/q*
$qO�/�/ �O�O�O�O�O__%_ 7_I_[_m__�_�_�_��_�? OOo5UM�P_OPTION �"./aTRW��&)�PePME��CoY�_TEMP  ?È�3B���`s�A�`�dUNI<��ŤaK�YN_BR�K U��t�EDITOR5a;a}o�b�_G@ENT 1V�N  ,&�PNS001.�A⤐ �E�&�MOVESAFE=�j3t5;�_3tc43��4s21� ��t��3u�)�3t#34D�V��t2p��� �to���g���ُ�uǏ ��u�1�3u�]��u�K���3t7w���&�APP_PALL�Oҟ�3s1�qB3LY���14'�9�����V�.EMGDI_STA�e���a� � +pNC�_INFO 1W<^�b���������ã��1X^� C��_8�+��
�do������ȿڿ� ���"�4�F�X�j�|� �Ϡϲ���������� ]e#�5�G�Y�g��g� �ߟ߱���������� �/�A�S�e�w��� ���������o��&� 8�J�\�v߀������� ��������"4F Xj|����� ���0BTn� x������� //,/>/P/b/t/�/ �/�/�/�/�/�/�/ (?:?L?f\?�?�?�? �?�?�?�? OO$O6O HOZOlO~O�O�O�O�O �O�O?? _2_D_�O p?z_�_�_�_�_�_�_ �_
oo.o@oRodovo �o�o�o�o�o�o�O_ *<Nh_r�� �������&� 8�J�\�n��������� ȏڏ��"�4�F� `j�|�������ğ֟ �����0�B�T�f� x���������ү��� ��,�>�X�J�t��� ������ο���� (�:�L�^�pςϔϦ� �����������$�6� P�b�l�~ߐߢߴ��� ������� �2�D�V� h�z����������  �
��.�@�Z�d�v� �������������� *<N`r�� ���F���& 8R�\n���� ����/"/4/F/ X/j/|/�/�/�/�/�/ ��/??0?JT?f? x?�?�?�?�?�?�?�? OO,O>OPObOtO�O �O�O�O�O�/�O__ (_B?8_^_p_�_�_�_ �_�_�_�_ oo$o6o HoZolo~o�o�o�o�o �O�O�o �oL_V hz������ �
��.�@�R�d�v� ���������o�o�� �*�DN�`�r����� ����̟ޟ���&� 8�J�\�n��������� ȯ�����"�<�F� X�j�|�������Ŀֿ �����0�B�T�f� xϊϜϮ���گ���� ��4�&�P�b�t߆� �ߪ߼��������� (�:�L�^�p���� �������� ��,�>� H�Z�l�~��������� ������ 2DV hz�������� �
6�@Rdv �������/ /*/</N/`/r/�/�/ �/"��/�/??. 8?J?\?n?�?�?�?�? �?�?�?�?O"O4OFO XOjO|O�O�O�O�/�O �O�O_&?0_B_T_f_ x_�_�_�_�_�_�_�_ oo,o>oPoboto�o �o�o�O�o�o�o_ :L^p��� ���� ��$�6� H�Z�l�~������o�o ؏�����(2�D�V� h�z�������ԟ� ��
��.�@�R�d�v� ������ƏЯ����  �*�<�N�`�r����� ����̿޿���&� 8�J�\�nπϒϤϾ� ���������"�4�F� X�j�|ߎߠ߲����� ������0�B�T�f� x������������ ��,�>�P�b�t��� ������������ (:L^p���� ������$6 HZl~���� ���/ /2/D/V/ h/z/�/���/�/�/ �/?.?@?R?d?v? �?�?�?�?�?�?�?O O*O<ONO`OrO�O�/ �/�O�O�O�O
?_&_ 8_J_\_n_�_�_�_�_ �_�_�_�_o"o4oFo Xojo|o�o�O�o�o�o �o_0BTf x������� ��,�>�P�b�t��� �o����Ώ���o��� (�:�L�^�p������� ��ʟܟ� ��$�6��H�Z�l�~��� �$�ENETMODE� 1Y��_�  �������ů׫��OAT�CFG Z���ܡ�ԢC���DATA 1�[����ա*F�*ݨd�v�����"��d��ʻ����ο ��
��.�@�R�d�޿ �ϬϾ�������n� ߒ�<�N�`�r߄ߖ� �"���������&� 8����n����� ��B���f��"�4�F� X�j�������������������RPOS/T_LO��]/����
�N`r���R�ROR_PR* �%��%����TA�BLE  ����	-RSE�V_NUM â?  ���]� _AUTO_ENB  ᥼��w_NOr ^���֡\  *�*�������h�+�����FLsTRz�HISY��񼠇_ALM �1_�� ������+��/�/�/��/�/�/�_R�  ���ע-:���TCP_VER �!��!��/$E{XT) _REQ.&s�3SIZ�?�z4STK�9���|2TOL  ���Dz6"�A z4_BWD0�0&�Aܢ�3DI�1 �`�9ء��KST�EP$O6O��P@OP�_DO�?��FAC�TORY_TUN�.'d�IDR_GR�P 1a��!d �	(?�Oנ�@�������gl�rw�q�����J ����V�C,_=]�@A��<B��%B���'AId�B��R@�"�B]@��s�B�=�B�H�@���A?��@!�l\�~=_@_�_�_vR��|�A0QA��S@�_�A�(\A*߰B]�����]�����ɡ��ul��8,4����B]<`�>�YBm@�I¡�~QBeBGc�_e"�Q�_��_�o�o�oHWC`}�dC��NqB�s{
uj^UUT&�UT�oO�o E׻� v�A^OH�cEP]��O���#M�˪qKA��B]?�p�d�:6:N���q9-��uB]���J��-p �1���<�����k;��FEATURE �b��@ۡ�Handlin?gTool e����Englis�h Dictio�naryk�4D ;StZ�arde�m��Analog I�/O����gle �Shift��ut�o Softwa�re Updat�e݉matic ?Backupi���ground E�dit^�k�Cam�era��F��Cn?rRndIm�G��ommon ca?lib UIB�j��n)�u�Monit�or��trc�Re�liab̀j�DH�CP^���ata ?Acquis����?iagnos���~ԛisplay,�?Licens�����ocument �Viewe����u�al Check Safety}�~n�hanced}�4j�o�sB�Fr:�l��xt. DIO 捐fi
���end.s�Err��L	���J��s��r���� �0�h�FCTN Me�nu[�v���TPw In��fac"�m�GigE4�F�"��p Mask Ekxco�g��HT2��Proxy Sv�C�}�igh-Spes�Ski]�~��~��mmunic�7ons��ur����ϟ��5�conne�ct 2�ncr4�stru����e9�S�J	�n�KA�REL Cmd.� Lx�uaz�I�R�un-Ti��Enyv?���el +
�s�S/Wk�$�V��B�РBook(S�ystem)h�M�ACROs,��/�OffseӀ��H0����͟��MR������MechStoEp��t����iˢ�ϋ>�xs������o}d̀witchl�����.�ƒ�Optqm��ӊ�filB���g���ulti�-Tp�,�i�PCMO fun��o�xV��:�Regi��Yrϰ�ri;�F*��r汀Num Se�l6Ս阠 Adj�u�����ϊ��ta�tun���=�m�RDM Robot|��scove���e�a���Freq �AnlyϷRem�4Э�n���&�Se�rvo���j�SN�PX b��ԎSN�2�Cli:���ЂLGibr����Z� E������o��t�ss#ag�n�A0 ����g�A0/I3�MI�LIB?P F�irm�)P�A�cc#�+�TPTXɟeln��\xb���*orqùimula��@��u��Pa��)"���:��&��ev.��riS��USB� port u�i�PĠa;�fR E�VNTYknexcepts�[�H�f,��y�VCy�rʲ��:�V��z�����S��SC�*/SG�E?/5%UIg�Web Pl��x.{����$��m�9��ZDT Applȴh��!EOAT%�l�y<�/7Grid*��\
=�/iR�.���^6����-200�0iC/125L~F�C-Link4��2�En�rk�n�l�x���Gu���?�2PT���s��tt���2���o;�e�E�yc�̀o�y�T`�-�maOin N��{�.
��RL���)~�MIo Dev%� (�� ��
�����`�/EB��Z�@t��miŠr�$�Ienp��G�4��asswoA3߁3���&n�64MB �DRAM�?xSFR9O�_7�ell��h�#sh�Q�_�Wc���U��p �\tỳs ��XLA�ЍB��Z�X��ҝ� 2%�a��<qn�MAIL�+l��@T���f�%�z�qf�T1����Д�VT?OPC-UA�s#T 2��O$QSĠn�Gcro��=�ṕ�yn.(RSS)�n���R4n��A�`ueCst��{P����S%Peˢtex�����;mi�Sp;�V��)PPs�à��i�dpnXy4�VRq�h� z�������ݏԏ��� 
�7�.�@�m�d�v��� ����ٟП����3� *�<�i�`�r������� կ̯ޯ��/�&�8� e�\�n�������ѿȿ ڿ���+�"�4�a�X� jϗώϠ��������� ��'��0�]�T�fߓ� �ߜ�����������#� �,�Y�P�b���� �����������(� U�L�^����������� ������$QH Z�~����� � MDV� z������/ 
//I/@/R//v/�/ �/�/�/�/�/??? E?<?N?{?r?�?�?�? �?�?�?OOOAO8O JOwOnO�O�O�O�O�O �O_�O_=_4_F_s_ j_|_�_�_�_�_�_o �_o9o0oBooofoxo �o�o�o�o�o�o�o 5,>kbt�� ������1�(� :�g�^�p��������� ʏ��� �-�$�6�c� Z�l���������Ɵ� ���)� �2�_�V�h� ��������¯���� %��.�[�R�d����� ����������!�� *�W�N�`ύτϖϨ� ����������&�S� J�\߉߀ߒߤ߶��� ������"�O�F�X� ��|���������� ���K�B�T���x� ������������ G>P}t�� ����C :Lyp���� ��	/ //?/6/H/ u/l/~/�/�/�/�/�/ ?�/?;?2?D?q?h? z?�?�?�?�?�?O�? 
O7O.O@OmOdOvO�O �O�O�O�O�O�O_3_ *_<_i_`_r_�_�_�_ �_�_�_�_o/o&o8o eo\ono�o�o�o�o�o �o�o�o+"4aX j|������ �'��0�]�T�f�x� ������������#� �,�Y�P�b�t����� ����������(� U�L�^�p��������� �ܯ���$�Q�H� Z�l�~��������ؿ ��� �M�D�V�h� zϧϞϰ�������� 
��I�@�R�d�vߣ� �߬���������� E�<�N�`�r���� ���������A�8� J�\�n����������������=, � H552�5[21aR78�`50aJ614�aATUP�54�5�6aVCAM�aCRI�UIFv�28�NREm�52�R63lS�CHaLIC�DwOCV!CSUm�869�0�EI�OC�4`R69��ESET��J�7�R68lMA{SKaPRXY�]7aOCO�3�h`��3�J6��53DH�LCH^�OPLG�0��MHCR�S?'MkCS�0�55��MDSW�'�OP��MPR�(0n�PCM�R0�'���I '51�5u1 80�PRS��69�FRD�FwREQmMCNa{93�SNBA�^�SHLBm6M�7t|(2�HTC��TMILmDTP�A\TPTX�6EL`6I D8wu lwJ95�TUT��95�UEV�U�EC�UFR�V�CChHOX&VIP��6CSC�6CSGt�6IaWEB�7HTT�R6�Hl� �FCG�GIG�GoIPGS�FRC�6�DG�H72�7�8�61�R53v�'68�R66��0��0�75�R65l55��P|Wk76�7l64 G�5�WR76�D0u6�F�XCLI�(��CMS\-`�S[TY�GTO�G7C�� |WNNli�ORSX&��M.8� 8�OPIVSEND��7`gLsGS�j7n�ETS�gLM088G�0�IPN�5< ?Qcu���� �����)�;�M� _�q���������ˏݏ ���%�7�I�[�m� �������ǟٟ��� �!�3�E�W�i�{��� ����ïկ����� /�A�S�e�w������� ��ѿ�����+�=� O�a�sυϗϩϻ��� ������'�9�K�]� o߁ߓߥ߷������� ���#�5�G�Y�k�}� ������������� �1�C�U�g�y����� ����������	- ?Qcu���� ���);M _q������ �//%/7/I/[/m/ /�/�/�/�/�/�/�/ ?!?3?E?W?i?{?�? �?�?�?�?�?�?OO /OAOSOeOwO�O�O�O �O�O�O�O__+_=_ O_a_s_�_�_�_�_�_ �_�_oo'o9oKo]o oo�o�o�o�o�o�o�o �o#5GYk} ����������1�C�  �H552E�_�2�1e�R78d�50�e�J614e�AT�UP��545��6�e�VCAMe�CR�I�UIF��28n�NREu�52ԊwR63t�SCHe��LIC$�DOCV�e�CSUu�869z��0��EIOC%��4d�R69ԊES�ET��ӋJ7ӋR{68t�MASKe��PRXY�7e�OCO�3��d�񐔌m3D�J6��53���H��LCH$�OP�LG��0d�MHCuR%�S�MCS���0��55��MDS�WE�S�OPS�MP�RT�A���0��PCM�R0��񐤊񠶔�51ċ51�0nĊPRS�69D��FRD�FREQnu�MCNe�93���SNBA5���SH�LBu�M��A�4�2HTC��TMI�Lu���TPA��T7PTX��ELd��┛8����t�J95n�TUTT�95D�wUEV�UEC$�wUFR�VCC���O�VIP��CS�C$�CSG$���I�e�WEB��HTT���R63�Rܱ�$�C�GC�IG#�IPGmS��RC��DGS��H72t�78��6�1�R53Ի68.��R66d�0���vd�75ĊR65t�c55d�q�4�76���7t�64d�5��R�76ĊD06��F���CLI��ËCMqS��! ��STY�ۋTOD�7��1�4�N9NtD�ORS��┊M"�q���OPI^��SEND5�7d�L��S�7D�ETS�LM$�C���$�IPN��D���� ����	//-/?/ Q/c/u/�/�/�/�/�/ �/�/??)?;?M?_? q?�?�?�?�?�?�?�? OO%O7OIO[OmOO �O�O�O�O�O�O�O_ !_3_E_W_i_{_�_�_ �_�_�_�_�_oo/o AoSoeowo�o�o�o�o �o�o�o+=O as������ ���'�9�K�]�o� ��������ɏۏ��� �#�5�G�Y�k�}��� ����şן����� 1�C�U�g�y������� ��ӯ���	��-�?� Q�c�u���������Ͽ ����)�;�M�_� qσϕϧϹ������� ��%�7�I�[�m�� �ߣߵ���������� !�3�E�W�i�{��� ������������/� A�S�e�w��������� ������+=O as������ �'9K]o �������� /#/5/G/Y/k/}/�/ �/�/�/�/�/�/?? 1?C?U?g?y?�?�?�? �?�?�?�?	OO-O?O QOcOuO�O�O�O�O�O �O�O__)_;_M___ q_�_�_�_�_�_�_�_ oo%o7oIo[omoo �o�o�o�o�o�o�o !3EWi{�� �������/��A�M�STD~H�LANGi� d�|�������ď֏� ����0�B�T�f�x� ��������ҟ���� �,�>�P�b�t����� ����ί����(� :�L�^�p��������� ʿܿ� ��$�6�H� Z�l�~ϐϢϴ�����p����� �RBTh�OPTN=�O�a�s߀�ߗߩ߻�����i�DPNg���'�9�K� ]�o��������� �����#�i�@�G�Y� k�}������������� ��1CUgy �������	 -?Qcu�� �����//)/ ;/M/_/q/�/�/�/�/ �/�/�/??%?7?I? [?m??�?�?�?�?�? �?�?O!O3OEOWOiO {O�O�O�O�O�O�O�O __/_A_S_e_w_�_ �_�_�_�_�_�_oo +o=oOoaoso�o�o�o �o�o�o�o'9 K]o����� ����#�5�G�Y� k�}�������ŏ׏� ����1�C�U�g�y� ��������ӟ���	� �-�?�Q�c�u����� ����ϯ����)� ;�M�_�q��������� ˿ݿ���%�7�I� [�m�ϑϣϵ����� �����!�3�E�W�i� {ߍߟ߱��������� ��/�A�S�e�w�� ������������ +�=�O�a�s������������������	�-?
99A�$�FEAT_ADD ?	���p�x   	 @������� �#5GYk} �������/ /1/C/U/g/y/�/�/ �/�/�/�/�/	??-? ??Q?c?u?�?�?�?�? �?�?�?OO)O;OMO _OqO�O�O�O�O�O�O �O__%_7_I_[_m_ _�_�_�_�_�_�_�_ o!o3oEoWoio{o�o �o�o�o�o�o�o /ASew��� ������+�=� O�a�s���������͏ ߏ���'�9�K�]� o���������ɟ۟� ���#�5�G�Y�k�}� ������ůׯ���� �1�C�U�g�y����� ����ӿ���	��-��?�Q�c�cDEMO� bp	   @�͠ϲ����� �����K�B�T�n� xߥߜ߮�������� ��G�>�P�j�t�� ������������ C�:�L�f�p������� ������	 ?6 Hbl����� ��;2D^ h������/ �
/7/./@/Z/d/�/ �/�/�/�/�/�/�/? 3?*?<?V?`?�?�?�? �?�?�?�?�?O/O&O 8ORO\O�O�O�O�O�O �O�O�O�O+_"_4_N_ X_�_|_�_�_�_�_�_ �_�_'oo0oJoTo�o xo�o�o�o�o�o�o�o #,FP}t� �������� (�B�L�y�p������� ���܏���$�>� H�u�l�~�������� ؟��� �:�D�q� h�z�������ݯԯ� �
��6�@�m�d�v� ������ٿп��� �2�<�i�`�rϟϖ� �����������.� 8�e�\�nߛߒߤ��� ��������*�4�a� X�j���������� ����&�0�]�T�f� ���������������� ",YPb�� ������ (UL^���� ���� //$/Q/ H/Z/�/~/�/�/�/�/ �/�/�/? ?M?D?V? �?z?�?�?�?�?�?�? �?OOIO@OROOvO �O�O�O�O�O�O�O_ _E_<_N_{_r_�_�_ �_�_�_�_�_
ooAo 8oJowono�o�o�o�o �o�o�o=4F sj|����� ���9�0�B�o�f� x�������ۏҏ��� �5�,�>�k�b�t��� ����ןΟ�����1� (�:�g�^�p������� ӯʯܯ�� �-�$�6� c�Z�l�������Ͽƿ ؿ���)� �2�_�V� hϕόϞ��������� ��%��.�[�R�dߑ� �ߚ��߾�������!� �*�W�N�`���� �����������&� S�J�\����������� ������"OF X�|����� �KBT� x������/ //G/>/P/}/t/�/ �/�/�/�/�/??? C?:?L?y?p?�?�?�? �?�?�?	O OO?O6O HOuOlO~O�O�O�O�O �O_�O_;_2_D_q_ h_z_�_�_�_�_�_o �_
o7o.o@omodovo �o�o�o�o�o�o�o 3*<i`r�� ������/�&� 8�e�\�n��������� ȏ�����+�"�4�a� X�j���������ğ� ���'��0�]�T�f� �������������� #��,�Y�P�b����� ����������� (�U�L�^ϋςϔϮ� ����������$�Q� H�Z߇�~ߐߪߴ��� ������ �M�D�V� ��z���������� �
��I�@�R��v� ������������ E<N{r�� ����A 8Jwn���� ��/�/=/4/F/ s/j/|/�/�/�/�/�/ ?�/?9?0?B?o?f? x?�?�?�?�?�?�?�?�O5O,O>OkObO�M  �H�O�O�O �O�O�O_"_4_F_X_ j_|_�_�_�_�_�_�_ �_oo0oBoTofoxo �o�o�o�o�o�o�o ,>Pbt�� �������(� :�L�^�p��������� ʏ܏� ��$�6�H� Z�l�~�������Ɵ؟ ���� �2�D�V�h� z�������¯ԯ��� 
��.�@�R�d�v��� ������п����� *�<�N�`�rτϖϨ� ����������&�8� J�\�n߀ߒߤ߶��� �������"�4�F�X� j�|���������� ����0�B�T�f�x� �������������� ,>Pbt�� �����( :L^p���� ��� //$/6/H/ Z/l/~/�/�/�/�/�/ �/�/? ?2?D?V?h? z?�?�?�?�?�?�?�? 
OO.O@OROdOvO�O �O�O�O�O�O�O__ *_<_N_`_r_�_�_�_ �_�_�_�_oo&o8o Jo\ono�o�o�o�o�o �o�o�o"4FX j|������ ���0�B�T�f�x� ��������ҏ���� �,�>�P�b�t����� ����Ο�����(� :�L�^�p��������� ʯܯ� ��$�6�H� Z�l�~�������ƿؿ ���� �2�D�V�h�|zό�  �� ���Ϻ��������� &�8�J�\�n߀ߒߤ� �����������"�4� F�X�j�|������ ��������0�B�T� f�x������������� ��,>Pbt ������� (:L^p�� ����� //$/ 6/H/Z/l/~/�/�/�/ �/�/�/�/? ?2?D? V?h?z?�?�?�?�?�? �?�?
OO.O@OROdO vO�O�O�O�O�O�O�O __*_<_N_`_r_�_ �_�_�_�_�_�_oo &o8oJo\ono�o�o�o �o�o�o�o�o"4 FXj|���� �����0�B�T� f�x���������ҏ� ����,�>�P�b�t� ��������Ο���� �(�:�L�^�p����� ����ʯܯ� ��$� 6�H�Z�l�~������� ƿؿ���� �2�D� V�h�zόϞϰ����� ����
��.�@�R�d� v߈ߚ߬߾������� ��*�<�N�`�r�� ������������ &�8�J�\�n������� ����������"4 FXj|���� ���0BT fx������ �//,/>/P/b/t/ �/�/�/�/�/�/�/? ?(?:?L?^?p?�?�? �?�?�?�?�? OO$O 6OHOZOlO~O�O�O�O �O�O�O�O_ _2_D_ V_h_z_�_�_�_�_�_ �_�_
oo.o@oRodo vo�o�o�o�o�o�o�o *<N`r� �������� &�8�J�\�n������� ��ȏڏ����"�4� F�X�j�|�������ğ ֟�����0�B�T� f�x���������ү� ����,�>�P�b�t� ��������ο��� �(�:�L�^�pςϑ����ȬϾ����� ����*�<�N�`�r� �ߖߨߺ�������� �&�8�J�\�n��� ������������"� 4�F�X�j�|������� ��������0B Tfx����� ��,>Pb t������� //(/:/L/^/p/�/ �/�/�/�/�/�/ ?? $?6?H?Z?l?~?�?�? �?�?�?�?�?O O2O DOVOhOzO�O�O�O�O �O�O�O
__._@_R_ d_v_�_�_�_�_�_�_ �_oo*o<oNo`oro �o�o�o�o�o�o�o &8J\n�� �������"� 4�F�X�j�|������� ď֏�����0�B� T�f�x���������ҟ �����,�>�P�b� t���������ί�� ��(�:�L�^�p��� ������ʿܿ� �� $�6�H�Z�l�~ϐϢ� ����������� �2� D�V�h�zߌߞ߰��� ������
��.�@�R� d�v��������� ����*�<�N�`�r� �������������� &8J\n�� ������" 4FXj|��� ����//0/B/ T/f/x/�/�/�/�/�/ �/�/??,?>?P?b? t?�?�?�?�?�?�?�? OO(O:OLO^OpO�O��I�$FEAT_�DEMOIN  ��D��@��@��DINDEX�K��A��@ILECO�MP c����A�B�E�@�SETUP2 �d�ER� � N /Q�C_AP2BCK 1e�I?  �)�Hc_"r[%Y_�_�@�@�_ �_�EX_�_|_o�_o Go�_ko�_�o�o0o�o To�o�o�o�oCU �oy�,��b ���-��Q��u� �����:�Ϗ�p�� ��)���6�_��� ����H�ݟl����� 7�Ɵ[�m����� ��� D�¯�z����3�E� ԯi�������.�ÿR� �����Ϭ�A�пN� w�ϛ�*Ͽ���`��� ���+ߺ�O���s߅� ߩ�8���\����� '��K�]��߁��� ��F���j������5����Y���f���	Y=PP�A_ 2VP*.cVR����N�*���	K�3���PC�;dN�FR6:DO��CT�@ ��y��@�:�*.F��kM�	{Y�'�KSTM��x~ �"-�@/KH/s/�'a//0/�/LGIF�/�/%�/�/�/I?LJPGS?}?%i?0&?8?�?D
JS�? O�N��3�?�?%
J�avaScript,OW?CSO�O&�qO.O %Cas�cading S�tyle She�ets�O"�
AR�GNAME.DT�OB� \�O�OA�#T4_�O#PDISP**_@�Tz_8_�JQ�Q�_d_
PANEL1/oS�_�_�QiPendant Panel<o"�	+d�_o'h�oDoVo�o�W21o%h �o�omxi2�o�@�h�J\��Y39�"�%h���u�xi3 ����h��R�d����Y4A�*�%h�֏�}�xi4ŏ���h��Z�l����DTPEINS�.XML�/�:\��ٟQCusto�m Toolba�r\�kYPASSW�ORD͟@�FR�S)a��`�Pas�sword Config��)��� "�_�u��������H� ݿl��Ϣ�7�ƿ[� ����� ϵ�DϮ��� z�ߞ�3�E���i��� �ߟ�.���R���v߈� ��A���:�w��� *����`�����+� ��O���s�����8� ��\�����'��K ]�����F� j���5�Y� R��B��x /�1/C/�g/��/ /,/�/P/�/t/�/? �/??�/c?u??�?(? �?�?^?�?�?O�?�? MO�?qO OjO�O6O�O ZO�O_�O%_�OI_[_ �O__�_2_D_�_h_ �_�_�_3o�_Wo�_{o �oo�o@o�o�ovo �o/�o�oe�o� ��N�r��� =��a�s����&��� J�\�񏀏����K��ڏo���$FIL�E_DGBCK �1e��b���� < ��)
SUMMA�RY.DG�+��MD:���7��Diag Sum�mary���
C?ONSLOG�̟�ޑ7�w�� �so�le lo���	?TPACCNm�ү�%�����TP �Accounti�n���FR6:�IPKDMP.ZIP+�/�
C�|����Excepti�on��1�ߐMEMCHECK�T������Memor?y Data�X��(i�)	FTAPj�[��_�����mment TB�D��8�s�T)�ETHERNET�}�)�±����E�thernet ~��figura����r�DCSVRF�|�b�tύ��%�R� verify� all��;ĸ�=�M�DIFF��k߸}���%��d�iff���±R�CHG01	����ﰢ�*����`�U�2 ��t���&����\��3���
��� �1���U�VTRNDIAG.LS���|���#��� O�pe3� Log ~�nostic8����<)VDEV��DAT$�%��VisFD�eviceMZIMG��r���),�=�Imag�X7UPp ESo?FRS:\o���Update?s List���FLEXEV�EN�3/���� UIF Ev��J 4/?�w�$)�
PSRBWLD'.CM_/+��w/����PS_ROB�OWEL��?�:GIGEJϐ//7?�GigEOY/<�7�x�M�SMHϕ?�$?�?��1/Em�ail��ae?s5��L)�1HADO�W�?�?�?AO�S�hadow Ch�angesDO;� ���BRCMERAR9OO0O�O��@�CFG Erro�r� t�0hO ������@SGLI�B�O�O�OK_N2U �St4�T�OQ��)7PZD�?�_4_��_�ZDI ad�k_�L~�)�PI�RDG_REPO�R��_�_�_%�iRPs Rep�or� ���BNOTIW�,o>o��o�Notif�ic4��_9���( �*1�NU�[�� �7��m��&� 8��\������!��� E�ڏi�����4�Ï X�j��������ğS� �w�����B�џf� ��s���+���O���� �����>�P�߯t�� ����9�ο]�򿁿�� (Ϸ�L�ۿpς�Ϧ� 5�����k� ߏ�$�6� ��Z���~�ߋߴ�C� ��g�����2���V� h��ߌ�����Q��� u�
����@���d��� ����)���M������� ��<N��r� %��[�& �J�n��3 ��i��"/�// X/�|//�/�/A/�/ e/�/?�/0?�/T?f? �/�??�?=?�?�?s? O�?,O>O�?bO�?�O �O'O�OKO�O�O�O_ �O:_�OG_p_�O�_#_ �_�_Y_�_}_o$o�_ Ho�_lo~oo�o1o�o Uo�o�o�o �oDV �oz	��?�c �
��.��R��_����i��$FILE�_FRSPRT � ��r�������MDONLY 1e��~i� 
 �� �A��e�%�N��r� �����7�̟[��� ��&���J�\�럀�� ��3���گi�����"� 4�ïX��|������ A�ֿ�w�ϛ�0Ͽ� =�f�����Ϯ���O� ��s��ߩ�>���b� t�ߘ�'߼�K�����~��VISBCKψ|��ރ*.VD��|C��FR:\��ION\DATA�\.�����Vi�sion VD fileo�}߷��� ���������"�G��� k������0���T��� x�����CUy �,��b�� -�Q�u �:���/�)/ �:/_/��//�/�/ H/�/l/?�/�/7?���LUI_CONF�IG f��|%�B; $  3Ԇ{���?�?�?�?�?�?I�0|x)?+O=O OOaOsO�LO�O�O�O �O�O�O�O$_6_H_Z_ l__�_�_�_�_�_�_ �_o o2oDoVoho�_ �o�o�o�o�o�o}o
 .@Rd�o�� ����y��*� <�N�`���������� ̏ޏu���&�8�J� �[���������ȟ_� ����"�4�F�ݟj� |�������į[���� ��0�B�ٯf�x��� ������W������ ,�>�տb�tφϘϪ� ��S�������(�:� ��^�p߂ߔߦ�=߷� ���� ��$��H�Z� l�~���9������� ��� ���D�V�h�z� ����5���������
 ��@Rdv�� 1����� <N`r��-� ���/�/8/J/ \/n/�//�/�/�/�/ �/�/�/"?4?F?X?j? |??�?�?�?�?�?�? �?O0OBOTOfOxOO �O�O�O�O�O�O�O_ ,_>_P_b_t__�_�_�_�_�_�_�X  �x�_c�$FL�UI_DATA �g���;a��Q-dRESULT 2h;e�d` �T��/wizard�/guided/�steps/Experto�o�o�o �o�o�o+=O�]z�Conti�nue with{ Gx`ance] ���������(�:�L�^� b-�a;e}�0 ���P}���;a�oops`������0�B� T�f�x�������mp�_ ՟�����/�A�S� e�w�������������t񯳌Ærip�` я7�I�[�m������ ��ǿٿ�����!�3� E�W�i�{ύϟϱ��� �������ʯܯ&�P��Ï�`Time?US/DSTߛ� �߿���������+��=�O�fwEnabl��������������%�7�I�[�by�3ߕ���i�{�24������!3 EWi{��^�p� ���/AS ew���l�~�������no�bditor�?/Q/c/u/�/�/��/�/�/�/�/b{ T�ouch Pan�el (# (re�commenz`) ?F?X?j?|?�?�?�?`�?�?�?�?i� ����=OOO/bacces+��O�O�O�O�O��O�O_"_4_F_a|�qpnect to� Network U_�_�_�_�_�_�_�_@
oo.o@oRoH��!QO3O�o��!gO% �IntroductionXo�o�o #5GYk}�� �������1��C�U�g�y���������oɏ���et�utojog!$Overview�� >�P�b�t��������� Ο����(�:�L� ^�p���������ʯܯ� � ��ӏ�G�r��"�$!SelmPT1Mod����� ��˿ݿ���%�7� I��m�ϑϣϵ��� �������!�3�E�� �(�rߜߺ�(c�$"~�TeachP/0antV�����&� 8�J�\�n����c� ���������"�4�F� X�j�|�����_ߡ߃�����l$��u�Join& g��@Rdv ��������� *<N`r�� �����������L5/G/�'!�r�`_'�/�/�/�/�/�/ �/??1?C?g?y? �?�?�?�?�?�?�?	O O-O?OQO/"/lO�O�X/n�HoldDe�admanSwitchRO�O�O_!_ 3_E_W_i_{_�_�_^? �_�_�_�_oo/oAo Soeowo�o�oZO�O~O��o�� �Ou�ResetAlarm�o 8J\n���� ����_�"�4�F� X�j�|�������ď֏�菧o�o�o�?�]�!8u�~%_J1���� ����ß՟����� /�A� �e�w������� ��ѯ�����+�=�N���i���g�?_J2-J6N�� ����,�>�P�b�t� �Ϙ�W���������� �(�:�L�^�p߂ߔ�`��e�w������#��Car�/3�E�W� i�{���������� ����/�A�S�e�w� ������������������:�C&�q*� ������� );��_q�� �����//%/�7/I/d/�/�CW�v_XJ/�/�/ �/?#?5?G?Y?k?}? �?N�?�?�?�?�?O O1OCOUOgOyO�O�O�\/n/�O�OT��/_Y-Z�O1_C_U_g_y_ �_�_�_�_�_�_�?	o o-o?oQocouo�o�o �o�o�o�o�O�O�O�8���*_Rotation�/��� ������)�;� �__�q���������ˏ ݏ���%�7��o`<��Tbon_ ۟����#�5�G�Y� k�}���N���ůׯ� ����1�C�U�g�y����J�\�n������� ���LastScreen��,�>� P�b�tφϘϪϼ��� �ϟ���(�:�L�^� p߂ߔߦ߸����ߛ� ����	�3��B��_�q� ������������ �%�7���[�m���� ������������!D3���9��!� �E����� (:L^p�A� ����� //$/ 6/H/Z/l/~/�/Oa s�/��/? ?2?D? V?h?z?�?�?�?�?�? ��?
OO.O@OROdO vO�O�O�O�O�O�O�/ _�/'_�/N_`_r_�_ �_�_�_�_�_�_oo &o8oI_\ono�o�o�o �o�o�o�o�o"4 �OU_y;_��� �����0�B�T� f�x���Io����ҏ� ����,�>�P�b�t� ��E��i˟���� �(�:�L�^�p����� ����ʯܯ�� ��$� 6�H�Z�l�~������� ƿؿ�������/�� V�h�zόϞϰ����� ����
��.��R�d� v߈ߚ߬߾������� ��*��3��W�� CϨ���������� &�8�J�\�n���?ߤ� ����������"4 FXj|;��_� ����0BT fx������� �//,/>/P/b/t/ �/�/�/�/�/��� �%?�L?^?p?�?�? �?�?�?�?�? OO$O �HOZOlO~O�O�O�O �O�O�O�O_ _2_�/ ??w_9?�_�_�_�_ �_�_
oo.o@oRodo vo5O�o�o�o�o�o�o *<N`r� C_U_g_��_��� &�8�J�\�n������� ��ȏ�oُ���"�4� F�X�j�|�������ğ ֟������B�T� f�x���������ү� ����,�=�P�b�t� ��������ο��� �(��I��m�/��� �ϸ������� ��$� 6�H�Z�l�~�=��ߴ� ��������� �2�D� V�h�z�9ϛ�]Ͽ�� ����
��.�@�R�d� v��������������� *<N`r� ��������� #��J\n��� �����/"/�� F/X/j/|/�/�/�/�/ �/�/�/??�' K?u?7�?�?�?�?�? �?OO,O>OPObOtO 3/�O�O�O�O�O�O_ _(_:_L_^_p_/?y? S?�_�_�?�_ oo$o 6oHoZolo~o�o�o�o �o�O�o�o 2D Vhz�����_ �_�_�_��_@�R�d� v���������Џ�� ���o<�N�`�r��� ������̟ޟ��� &���	�k�-����� ��ȯگ����"�4� F�X�j�)�������Ŀ ֿ�����0�B�T� f�x�7�I�[������ ����,�>�P�b�t� �ߘߪ߼�{������ �(�:�L�^�p��� ������������ 6�H�Z�l�~������� �������� 1�D Vhz����� ��
��=��a #�������� //*/</N/`/r/1 �/�/�/�/�/�/?? &?8?J?\?n?-�?Q �?uw?�?�?O"O4O FOXOjO|O�O�O�O�O �/�O�O__0_B_T_ f_x_�_�_�_�_?�_ �?oo�O>oPoboto �o�o�o�o�o�o�o �O:L^p�� ����� ���_ o�_?�i�+o������ Ə؏���� �2�D� V�h�'������ԟ ���
��.�@�R�d� #�m�G�����}���� ��*�<�N�`�r��� ������y�޿��� &�8�J�\�nπϒϤ� ��u��������ϯ4� F�X�j�|ߎߠ߲��� �������˿0�B�T� f�x���������� ����������_�!� �������������� (:L^�� ����� $ 6HZl+�=�O�� s����/ /2/D/ V/h/z/�/�/�/o�/ �/�/
??.?@?R?d? v?�?�?�?�?}�?� O�*O<ONO`OrO�O �O�O�O�O�O�O__ %O8_J_\_n_�_�_�_ �_�_�_�_�_o�?1o �?UoO|o�o�o�o�o �o�o�o0BT f%_������ ���,�>�P�b�!o ��Eo��iok����� �(�:�L�^�p����� ����wܟ� ��$� 6�H�Z�l�~������� s�կ�����ϟ2�D� V�h�z�������¿Կ ���
�ɟ.�@�R�d� vψϚϬϾ������� �ů��3�]���� �ߨߺ��������� &�8�J�\�π��� �����������"�4� F�X��a�;߅���q� ������0BT fx���m��� �,>Pbt ���i�{�����/ ��(/:/L/^/p/�/�/ �/�/�/�/�/ ?�$? 6?H?Z?l?~?�?�?�? �?�?�?�?O��� SO/zO�O�O�O�O�O �O�O
__._@_R_? v_�_�_�_�_�_�_�_ oo*o<oNo`oO1O CO�ogO�o�o�o &8J\n��� c_�����"�4� F�X�j�|�������qo ӏ�o���o�0�B�T� f�x���������ҟ� ����,�>�P�b�t� ��������ί��� Ï%��I��p����� ����ʿܿ� ��$� 6�H�Z��~ϐϢϴ� ��������� �2�D� V��w�9���]�_��� ����
��.�@�R�d� v����k������� ��*�<�N�`�r��� ����g����������� &8J\n��� �������"4 FXj|���� �������'/Q/ x/�/�/�/�/�/�/ �/??,?>?P?t? �?�?�?�?�?�?�?O O(O:OLO/U///yO �Oe/�O�O�O __$_ 6_H_Z_l_~_�_�_a? �_�_�_�_o o2oDo Vohozo�o�o]OoO�O �O�o�O.@Rd v������� �_�*�<�N�`�r��� ������̏ޏ����o �o�oG�	n������� ��ȟڟ����"�4� F��j�|�������į ֯�����0�B�T� �%�7���[���ҿ� ����,�>�P�b�t� �Ϙ�W���������� �(�:�L�^�p߂ߔ� ��e��߉��߭��$� 6�H�Z�l�~���� ��������� �2�D� V�h�z����������� ��������=��d v������� *<N�r� ������// &/8/J/	k/-�/Q S/�/�/�/�/?"?4? F?X?j?|?�?�?_�? �?�?�?OO0OBOTO fOxO�O�O[/�O/�O �O�?_,_>_P_b_t_ �_�_�_�_�_�_�_�? o(o:oLo^opo�o�o �o�o�o�o�o�O�O�O E_l~��� ����� �2�D� oh�z�������ԏ ���
��.�@��oI #m���Y��П��� ��*�<�N�`�r��� ��U���̯ޯ��� &�8�J�\�n�����Q� c�u���鿫��"�4� F�X�j�|ώϠϲ��� ���ϧ���0�B�T� f�xߊߜ߮������� �ߵ�ǿٿ;���b�t� ������������ �(�:���^�p����� ���������� $ 6H��+�O� ���� 2D Vhz�K���� ��
//./@/R/d/ v/�/�/Y�/}�/� ??*?<?N?`?r?�? �?�?�?�?�?�??O &O8OJO\OnO�O�O�O �O�O�O�O�/_�/1_ �/X_j_|_�_�_�_�_ �_�_�_oo0oBoO foxo�o�o�o�o�o�o �o,>�O_!_ �E_G����� �(�:�L�^�p����� So��ʏ܏� ��$� 6�H�Z�l�~���O�� s՟矫�� �2�D� V�h�z�������¯ԯ 毥�
��.�@�R�d� v���������п⿡� �ş�9���`�rτ� �ϨϺ��������� &�8���\�n߀ߒߤ� �����������"�4� �=��a��Mϲ��� ��������0�B�T� f�x���I߮������� ��,>Pbt �E�W�i�{���� (:L^p�� ������ //$/ 6/H/Z/l/~/�/�/�/ �/�/�/���/?� V?h?z?�?�?�?�?�? �?�?
OO.O�ROdO vO�O�O�O�O�O�O�O __*_<_�/??�_ C?�_�_�_�_�_oo &o8oJo\ono�o?O�o �o�o�o�o�o"4 FXj|�M_�q_ ��_���0�B�T� f�x���������ҏ� ���,�>�P�b�t� ��������Ο���� �%��L�^�p����� ����ʯܯ� ��$� 6���Z�l�~������� ƿؿ���� �2�� S��w�9�;ϰ����� ����
��.�@�R�d� v߈�G��߾������� ��*�<�N�`�r�� Cϥ�g�������� &�8�J�\�n������� ����������"4 FXj|���� ������-��T fx������ �//,/��P/b/t/ �/�/�/�/�/�/�/? ?(?�1U??A �?�?�?�?�? OO$O 6OHOZOlO~O=/�O�O �O�O�O�O_ _2_D_ V_h_z_9?K?]?o?�_ �?�_
oo.o@oRodo vo�o�o�o�o�o�O�o *<N`r� ������_�_�_ #��_J�\�n������� ��ȏڏ����"��o F�X�j�|�������ğ ֟�����0��� �u�7�������ү� ����,�>�P�b�t� 3�������ο��� �(�:�L�^�pς�A� ��e��ω��� ��$� 6�H�Z�l�~ߐߢߴ� ��������� �2�D� V�h�z�������� ��������@�R�d� v��������������� *��N`r� ������ &��G	�k-�/� �����/"/4/ F/X/j/|/;�/�/�/ �/�/�/??0?B?T? f?x?7�?[�?�?�/ �?OO,O>OPObOtO �O�O�O�O�O�/�O_ _(_:_L_^_p_�_�_ �_�_�_�?�?�?�_!o �?HoZolo~o�o�o�o �o�o�o�o �OD Vhz����� ��
���_%o�_I� s�5o������Џ�� ��*�<�N�`�r�1 ������̟ޟ��� &�8�J�\�n�-�?�Q� c�ů������"�4� F�X�j�|�������Ŀ �������0�B�T� f�xϊϜϮ����ϑ� �����ٯ>�P�b�t� �ߘߪ߼�������� �տ:�L�^�p��� ��������� ��$� �����i�+ߐ����� �������� 2D Vh'�y���� ��
.@Rd v5��Y��}��� //*/</N/`/r/�/ �/�/�/�/��/?? &?8?J?\?n?�?�?�? �?�?��?�O�4O FOXOjO|O�O�O�O�O �O�O�O__�/B_T_ f_x_�_�_�_�_�_�_ �_oo�?;o�?_o!O #o�o�o�o�o�o�o (:L^p/_� ����� ��$� 6�H�Z�l�+o��Oo�� Ï����� �2�D� V�h�z�������� ���
��.�@�R�d� v���������}�Ǐ�� ��׏<�N�`�r��� ������̿޿��� ӟ8�J�\�nπϒϤ� �����������ϯ� �=�g�)��ߠ߲��� ��������0�B�T� f�%ϊ��������� ����,�>�P�b�!� 3�E�W߹�{����� (:L^p�� ��w��� $ 6HZl~��� �������/��2/D/ V/h/z/�/�/�/�/�/ �/�/
?�.?@?R?d? v?�?�?�?�?�?�?�? OO���]O/�O �O�O�O�O�O�O__ &_8_J_\_?m_�_�_ �_�_�_�_�_o"o4o FoXojo)O�oMO�oqO �o�o�o0BT fx�����o� ���,�>�P�b�t� ��������{oݏ�o� �o(�:�L�^�p����� ����ʟܟ� ��� 6�H�Z�l�~������� Ưد����͏/�� S���������¿Կ ���
��.�@�R�d� #��ϚϬϾ������� ��*�<�N�`���� C��߷�{������� &�8�J�\�n���� ��u��������"�4� F�X�j�|�������q� �ߕ���	��0BT fx������ ���,>Pbt �������/ ����1/[/�/�/ �/�/�/�/�/ ??$? 6?H?Z?~?�?�?�? �?�?�?�?O O2ODO VO/'/9/K/�Oo/�O �O�O
__._@_R_d_ v_�_�_�_k?�_�_�_ oo*o<oNo`oro�o �o�o�oyO�O�O�o�O &8J\n��� ������_"�4� F�X�j�|�������ď ֏�����o�o�oQ� x���������ҟ� ����,�>�P��a� ��������ί��� �(�:�L�^���A� ��e�ʿܿ� ��$� 6�H�Z�l�~ϐϢϴ� ſ������� �2�D� V�h�zߌߞ߰�o��� ���߷��.�@�R�d� v����������� ���*�<�N�`�r��� ���������������#��GY�$FM�R2_GRP 1�iY� ��C4  B]��	 ����� E�� ���� OHcEP]���O��#M{���KA����?� � :�6:N�;9-��C�A�  �_qBH�C`}�dC��N�B�{����ޔ @UUT�UT���/�>FD��>�d�>D��=�=��1�/5�H$:���=:��:.��	:sf�:�Uf��/C/}/�/�/�/��/�/�m_CFG� jzT �	?J?\?n?;NO �z

E157785   <�RM_CHKTYP  j�� � �Z lROM�0_MsIN�0����0u��Xm SSB 3�kY �O�C>OPO5�TP_DEF_O/W  ��eG�IRCOM�0vO��$GENOVRD�_DO�6�MT[HR�6 d�Ed�Do_ENB�O �@�RAVCslG�@ ���� ��}EӤ�G
��F�/lGC�,�/:Ok_�� #�0�E�q_���R�	QOUv r�z�1�zB�<�0!�_�_�_o,Co�C�i`�Yo�XL�o�lBȁo�a�cp�	�YWO
PSMTs�sY� @hd�$HoOSTC 21tz	n@�� 	>xM>{>�n�e����� �z�"�4�F�X�{|���	anonymous�����я��� =Oa>�u�� ������������� ��(�K�����p��� ���������#�5�7� $�k�H�Z�l�~���ן ��ƿؿ����U�g� D�V�h�zό�ӯ��� �����?��.�@�R� ��c߈ߚ߬߾����� )���*�<�N�ϧ� �����ߧ������� �&�m�J�\�n����� ������������" i�{��;����� �����0B Twx������ �+=Oa>/u� t/�/�/�/�/�/�/ ??(?K/��p?�? �?�?�?�/#/5/7? $Ok/HOZOlO~O�O�/ �O�O�O�OO�OU?2_�D_V_h_z_�o qEN�T 1u�[ P�!_�_  �`��P92.168.115.231�_ �_o�X8o�_\ono 1o�oUo�oyo�o�o�o �o�o4�oX|? �cu����� �B��;�)�g���_� ����䏧��ˏ,�>� �b�%���I���m�Ο �����ǟ(��L���p�3�E��� !Q�UICC0����!1�Z7ϯ���_ӯ��F���2H�$�6����!ROUTER�t����!PC�JOG�ÿ!��0.10����C�AMPRT8��!a�1�_�F�RT���c�u��� !So�ftware O�perator Panel��%�&���TNAME !��Z!
ROBOT�rac2��ZS_�CFG 1t�Y� �Au�to-start{ed�4FTP�?��O_��7O� � 2�D�V�Oz���� ����g���
��.�@� �>�ߪ߼ߙ����߰� ������;M_ q���(���� �?�?�?�?� ��������/ !/3/E/W/z��/�/ �/�/�/�/.@R/? f/S?�w?�?�?�?t/ �?�?�?OO<?�?8O aOsO�O�O�O�/?? &?(O_\?9_K_]_o_ �_HO�_�_�_�_�__ �_#o5oGoYoko}o�O �O�O�o�_�o0_ 1C
o y��� �o�f�	��-�?� �o�o�o�o����oϏ �����;�M�_� q�����(���˟ݟ� ��Z�l�~�,���� Ə����ǯٯ믲�� !�3�E�h�i�������౿ÿտi�=�_ER�R vG����P�DUSIZ  jv�^����>%�?WRD ?��W���  guestv�e�wω��ϭϿ�6�SCDMNGRP 2w��w��W�Tv�p�/v�0v�K�� 	P01.0�0 8<�   �A  %  �
��8�}=���2� �����������h`�}1`Ѓ���XL��  �8�� � �I��L��y�`��E���R����t��8�����=���
�=�V���{`���-p�Ռd�ep�����J$��B��$��d0��B�T�f���_GROUU��x�����	��'Ә�QUPD'  S������TY{����T�TP_AUTH �1y� <!iPendan���A���O� !KAREL:*A�J�\�KCq������i�VISION SET������v�g��� f�D2 \V�z������CTRL z���*
v�F�FF9E3�U��FRS:DEFA�ULTOFA�NUC Web ?ServerO= ����M�_�������//�WR_�CONFIG �{�� uO��I�DL_CPU_P5Cnv�B�X�� � B�9cy#MI�N�,=� ?�y~y GNR_IO���3�v�
�y NPT_�SIM_DO�&��+STAL_SC�RN�& ��*TPMODNTOL	7�+�RTY�(�!�&����ENB	7���u$OLNK 1|�a��?�?�?�?�?��?O}2MASTE�� ��}2SLAVE� }�4ERAM�CACHE#O��I}O�O_CFGeO�wIUO���OyBCMT_OPn�"ʻC�YCLdO�Eh_A�SG 1~��?�
 O*_<_N_`_r_ �_�_�_�_�_�_�_o�oK�BNUM2���
yBIPbOtGR?TRY_CN�O�EP1��2Ø1�� yB�@�BCNY��oY��y RCA_ACC� 2���  V�vq��j � � �� 6� W6�hv�'v�v��vZ 2�b�	u	�v�8|�dB�UF001 2����= l`u1�  u1l��t��u2�p2l��tಊsm�p�r uIuW3m@�sm�tm�t�m��t��t��snV�tn �t@�t`�tV�tn��sn�tn�tUo�to�to�o	�_p t� Q�p�t5p�tp�tp�J��tUp�tp�tq�tq�tUq�q�tqq�q�toq�p)�pi�t�i�u3F�.Q�j�p/�E�j ��sj�tj�tj�tj*�tj�tj�tk�p�qUk�tk�k�tk�tUk�tk�tk�tl�t%l�l�gy2t� �������� (�:�L�^�p��������C�1����qA����ЁÑ؁������ʐ�qZ���hA��
��.�@��R�d�ms3}���  ���������������  ������ʒ�����ٓ���������  �� �� �
� ��� ���!� ���1�   9�@��I�@��Y�`� �i�`���y�`�봉� `�������ĩ����� �������נ�ЁB� ؁�������ߠ ���ߠ��!�(��1� (Л�A�(��Q�(����a�����q�ev�A2����4���B�B�<�B��оҿ��"�dHIuSqr��� �q� 2023-0�3-2��B� P�2���"��� �Q(����8�@�AH���Џ��`��:q��À 9 q��; y2���<���Vu�`�؝� 	��-�?�Q�c�u��Ux��������U���������e���E��Vt�� �����	��-�?�Q�� * e� �1 m� 7 �u�����%ps��19��������) _�q�_q��r�
� ������	P-?Q%pq�
7u �������/(/)/��p�
6Q/c/ u/�/�/�/�/�/�/�/ ?����|�����/?A?�S?e?w?�?s� . ��L��O�O�O ��,O>OPObOtO�O�? �?�?�?�?����_(_�:_L_^_p_�P � 1A %  >$�P��d�P���_�_ }��_�_o o2oDo z_�_�_�oUg�o�o �o�o
.@Rd v?/������ ��*�<�N�?)?�� ������̏ޏ�����&��?�х�OOT�	UmR�\�\� \�U(\�0\�8\�@\�UH\�P\�X\�`\�=h\�p 	���ţ ү�����OQ�c�u����������:�x8���8��8��8��8���8��8��8��8��`9��_-�.;��G� �O��W��_��g� �o��w���� �»��à§�O��d��ſ׿鼯o 
��.�@�R�d�v��� �������£��� ���³��»������ ������	��-� ?�Q�c�u߇ߙ��g� ��������
��.�@� R�d�v��C������ ������
��.�@�R��R��4I_CFG �2�.� H
�Cycle Ti�meR�Bus}y�Idln^}min	���UpjpR�eadxDoYw�� �e�Countp	N'um e~�	��R���1PROG�K�.�8�� $i{�����	�R��0SDT_IS�OLC  .���  ��$J2�3_DSP_EN�B  �2� INC ��R� �Av�?֐=����<#�
!b):�o m!�/�/R��/,�/'OB?C$#f���M&�!G_GRO�UP 1��>qb< �b!(�&?�/?�Xe?R�Q{?�?�?�?�?�?��?OO��/�)G_IN_AUT���f�I* POSRE��/�&KANJI_�MASK�FlJKA�RELMON �.�R�y�?�O_@ _2_D_GN�BC�J�P"�fU�O�ECwL_L\@NUM( ��]�@EYLOGOGINGd�3��ra�M%:LANGUA_GE .�`��DEFAUgLT a�LGL��J� U������R��'�  � 
��R��R���;���
�a(UT13:\T_�o �o�o �o�o�o�o4ASe|R�(�O����PN_DISP ��E/�z?x??L�OCTOL�R�D�z4!^!'�GBOOK �!m���q��q�q����rh�� ������ˏ݋�-c���ۆ	E�pi"1��K�hnC�_BUF�F 2�� 	Y�N���^���� �Ɵ؟����;�2� D�q�h�z�������¯�ԯ���
�7��tADCS �JQ"f! ��;��8R����ÿտ�N�IO 2�Z�C W 
�W 4�� �0�B�V�f�xϊϞ� ������������.� >�P�b�v߆ߘߪ߾�~�ER_ITM�d<O�)�;�M�_�q� ������������ �%�7�I�[�m��!�N��SEV�@�}��TYP������8��}ARST�_L��SCRN_FL +2���4���������T�P�P����NG�NAM$$x�b�tU�PS�pGI4 �U�M%Z_LOAD�� G %%�ATTAUGHT�z@��MAXUA�LRM�R�A��rM%
�`_PRe��@ 9����C�p��!ot�����# 0Pw 2�O� ؞��	'��@ڤ@# ��tr"�/�/�/�/%( �/?�/'?
??]?H? �?l?�?�?�?�?�?�? �?�?5O OYODO}O�O rO�O�O�O�O�O_�O 1__U_g_J_�_v_�_ �_�_�_�_	o�_-o?o "ocoNo�ojo|o�o�o �o�o�o;&_ BT������ ���7��,�m�X� ��|���Ǐ���֏���DBGDEF ��
%!!�*�_LDXDISAE��MEMO_A�P?E ?
 <����������Ο������FR�Q_CFG ��
'@�A ��@�4]���<$d%����*�<�R"�
+^m$*Π/Т **:٢��̯ި w�����C�:�L�y� p�������
%ؿ��ɿ0���"��,(��V� ��Dρ�hϥό϶��� ������#�5��Y�@��}ߏ�v߳ߵISCg 1��� �� ��m$A����J�5�n������_MSTR ������SCD 1����f���b�� ��(��L�7�I���m� ��������������$ H3lW�{� �����2 VAf�w��� ���///R/=/ v/a/�/�/�/�/�/�/ �/??<?'?`?K?�? o?�?�?�?�?�?O�? &OO6O\OGO�OkO�O`�O�O�O�O��MK?�����q��O$MLoTARM>��E�)R �:�h_|pT)�METPUc���B����NDSP_ADCOL�U�o��^CMNT�_ ��UFN�P�_�WF�STLI�_�W�� ���?n_Sq�Woad��UPOSCFg��^PRPM�_qiS�T�P1��� 4i�#�
�a��e�o �g�o�o�oO1C �gy�������'�	��]�G��QS�ING_CHK � �_$MODAF=����'[)Y���DEV 	f�	�MC:�皂HS�IZEc��@ȗ�T�ASK %f�%�$1234567�89 8�J���TR�IG 1��� l)�v�������ǟ��F�YP��������EM_INF 1����`)AT&FV0E0̟�C�)+�E0V1�&A3&B1&D�2&S0&C1S�0=2�)ATZC���~�H��ïR����z�A��֯?�&�c�u� )���M�_�q� �������O�<�N�� r�-ϖϨϏ������ ߵ�ǿٿJ�U�π� �Ϥ�_�i��ߕ����� "�4���X���/�A� ��e���������0� ��T�f�M���=�O��� s�����>u� b'��S��� �����������p #����}����$//H/^ONIwTOR(`G ?ߋ�   	EX�EC1�C�"2�(3��(4�(5�([��&7*�(8�(9�C�" �$�"�$�"�$�"�$�" �$�"�$�"�$�"�$�"��$�"�#2�(2	82�82!82-82982�E82Q82]82i83��(3	83�"��R_�GRP_SV 1ݢ� (O�@�
s�z4 >���Q6tT��?�t?��]-"��_D��QCION�_DB������A�  ��@n�@o�&T�Dm`�Gɸ�@> ��> N �  ��@��L��m`>!)R-ud1��__+_�QPL_NAME !)��TP�!Def�ault Per�sonality� (from FsD)�@�RRR2A� 1�����$TQm`\ dRb�_�_�_�_�_�_ oo1oCoUogoyo�o �o�o�o�o�o�o	��2�_FXj|�@������B5 �$�6�H�Z�l�~��� ����Ə؏���� � 2�D�V�h�z������� ԟ���
��.�@� R�d�v���������Я �����*�<�N�`� r���������̿޿���&�5P<�N�`� rτϖϨϺ�����������}5P�@��\  �  ���  ��  A_�  BQ�TQЕ�5P
=АAБ���  ��@AL�B�Q�zQ��  C�5PC5PP E�;� E@ D����$�D|З՗�8|Уް��  �Փ�F��E�������g���E(�������Z���ӑ������$�/ �3�@�P���� � � p�����L������ќ�Ќ���P������������� � �������������P���@� �m��N�� �� ���l�� �����������	�P����������ЋҘ���$��$J�ᡢ�����H���a z|z�`�|�vFp E��0����FA3����2��B9����E��zE��ą5T*A  P�u�5Rdo9Ф ����X2Z��5WW%$�/N/&amB'l/b*ApM�=�u#����/i/T�/�' ��$Bh�@�.+@g@?<5RA%�	`V/P?b?t?31:�oAxR�?�?�?�>� �@�2h��&�X�A�D�A�@D3/� �5P�  ��5P� �� J��8�B7/XOCO|O�gOyO�O�O�O1^RR҃S�LY@@>2l�6 .2��� @��?|L�4Q��?��<4Q��@�6/�0�b^;�	lDR	�  <P� �,^@@}P��� � s? � � ��Rp�K�l,K����K��2KI+��KG0�K �U��Lb_�E��^�P@�6@ t�@�X@I� b�MP�_3�N�����
��ՙ�����`Pa�]��9eИ ��k���e���xa�_  �X�ￒ4������0o�Bxоo��Н��c':I>O�S��_q�$v�OB�E	'� � `r�I� �  ���!�J:�È~�È=��͜u�R@��p�nQ����R�<�o�JN<�0.�  'D�aE`?�� bQ`b�YoCm`BH�C4D��y`B�Ј������}����R� �P�� &�^;̀�HB� ܆�5�=�0 �q����O)��OM�8�0q�\�n�au5�rp������� ,��:�����Q
@�b�?��ff������ -0)�;��Q8��Q�_�K?�"�@Qd�(����P�����Q�S�T�s�|�����Q;�x5�;��0;�i�;�du;�t�<!���_��BT�SDR�0?fff�?�p?&>�4@׿�A#T�@�o[\��٨�9��� �P4U��2W��"�xT� �ӿ���0��T�?��xϊ�uϮϣر�F �0���ϙ�߅�/ߩ�h�b���E* C������<Q߲ߝ����� �����	��T�?�x� �?���i�__%���I� ���6�H�Z�l���� ��-������������1A�6� �"H�Am����?�؛���h�����s�W�C�>��` Ca���B��� �X `�l����bC@_;C�Ln�BA��Q�>V���������Y���\���
;�3��Q��hQ��@�G�B=ן
?h�ô� ���W�������B/
=�࿣��Ɗ=�K��=�J6XL�I�H�Y
H}��A�1��L�jL�LPBhH:���HK�,/> 	b�L �2J���H��H+UZBu��/� �/�/�/�/�/?�/3? ?C?i?T?�?x?�?�? �?�?�?�?�?/OOSO >OwObO�O�O�O�O�O �O�O__=_(_a_L_ ^_�_�_�_�_�_�_o �_o9o$o]oHo�olo �o�o�o�o�o�o�o# G2kV{�����yGϭ�� �C�aE� Ĉ��"�CVF��C�J��+��� ��K����� 
E�������	�� (��g_�h�ġ��<��u�N��,�>�j��3lC�X�j�x���ⷄ����t�.�3��}��k����q'�3�JJܝܙ�
�@�.�d��R��P��P��� �￯�˯��������&�_�J�o�{xo�~���  fU�� Z��ο��+�ү��0^�Lς�p�ψϒϘ�϶���)Z���� ? ( 5�9 ߀ �N�<�r�`ߖ߀� ? 2 E��Q�E�L�����q�QB�B 5�C�:*Y  @�
� Q ��)�;�M� �q���܌}��Ӥ`���������?��㈊���7�Q #���
 ��Q�c� u����������������);�������V{H��$M�R_CABLE �2��� 5Ȱ�T��@�?����� ' ´�л C� ���O4>�B������������I-C�{�5�����,  �����(��l��N�/�HB��-ܑw�ha 7�Hð�D3�jD��<�`���
�����B���&���B  "��;C��BG ���ԑ ��W��� ���C/>//`/8/ J/�/n/�/�/�/�/�/ �/??:??\?ړ"����� B���E�?�=ݏB�܍d�?�e�3�7�1������`��� �Ѡ���@�������� ����0��0��0����@�	������ ��0�	@��@� 2936/11  *MH} tOM ��	���'� ��<�i�(%% �2345678901�O�E ~O�O�A���������1���
�Gx=not� sentLK�C�W��TEST�FECSALGRO  eg~���dFTd��A
VT��謠�k���q_�_�_�_ �9UD1:\m�aintenan?ces.xm�_;� � '�]�DEFAUL�Ty�tGRP 2��eJ  �  ������ � �%!1st �cleaning� of cont�. vPilat�ion 56�R�B�cG�a�o��+s�����o�o�o}[d%�lamechs`c�al checkN`�Vs�`qg���o�����+v|aroller>Pb�k�X�j��|����+qBas�ic quarterly��'��j,G��&�8�J�\�#ycM5����"8��!�଑������� ���(�w�C�R���v��fϟ����ȯ�گ�+rGreas�e bal�Qr bush�f�;�����h�z�������+r�C�ge3r.
�t:y��  3"`�!��������	W�,��>�P�b�t�+qJ1� i-g�~�ge xϯ���"������&�8߇�2��c�u߇���#�ϴ��������߂��3R�'�9�K���$���x�����ﳂJ4/J5��� ���R(g�<�N�`�r������6��������U' +� $6H��Ⱥ�cabl���R�� �_��Re
��� ���ù|cտ��l���������Overh�au��c�" !x�P!/RewL/ ^/p/�/�/c�/�/�3 �)�/�X;/?"?4?F? X?�/|?�/�/�/�?�? �?�?OOm?BO�?�? �?�O�O�O�O�O!O�O _WO�O{OP_b_t_�_ �_�O�_�__�_A_o (o:oLo^o�_�o�_�_ �oo�o�o $so H�o�o~�o��� ��9�]oD�� h�z��������ԏ#� 5�
�Y�.�@�R�d�v� ŏ�����П���� �*�<���`�����ӟ ����̯ޯ��Q�&� u�����n��������� �m��;�ۿ_�4�F� X�j�|�˿�ϲ���� %�����0�Bߑ�f� ���Ϝ����������� �W�,�{ߍ�b�߆����� �/|��b 	 X=,�1?�V? ���=i�=�,����9X<7��4��>��B�(�B�qn<����>�;�A��  B�ff?@����B   =���?��#?�V>D�>�]d��T�<��S��-��>S�B��KC�s=�Hz?R;�s.�Rn�:�L�����?���>���>i�>�D���Q�:�o<�?���?�p�B|�n�B�G>[���@pbN.�S@O｢��>��%�?u>��7���,q�$��?	c>�M�=��2A7��B���>�$_�A<C�.��R��N>�<j?g�?^5?���333�i^�=��w>��>����"A	�B�ł6	��D��>����?^��R?���bE��<��Z>s��>���"��B�o����J� )�� i{ 6�Z�����O �Y�a@�� KGuaK�H!KH��K�Io�KJaK�J�!KKi�K�L�KL�aK�MnQKN K�N��KOl�K�P@KP� K�QkAKRK�E{!KF#�K�F̡!������`�� ��Ѡ��@�������� ��y ��} �� ����@�	����� ��y �� �� � �2026/1�1 *�) F�@ /$/6/H/Z/l/~/ �/�/�/�'m��/�/? ?&?8?J?\?n?�?�? �?�?�?�?�?�?O"O 4OFOXOjO|Cz�I� s_�_�_�__�_�_�_��}�yO�Fv�K�HQKH�K�Ip�KJ�K�J�QKKkK�L�KL��K�Mo�KNCK�N�KOm�K�P�KP�CK�Ql�KRDK�E|QKF%KF���O�O__*_�<_NR  ;�����$MR_HI_ST 2�V�p�� 
 \�$!1st c�leaning �of cont.� ventilation 56�`����ß��T�ǮG�V -3�19.4 hou�rs RUN 9��pqme�ch$pcal c�hecko�)� �m�"UK}�Oy950.3`x�vuu-qroll�er�����pBasic �quarterly����"�� �_Ώ������(�ߏ L�^����9�����o� ɟ�� ��$�۟�Z��l�~�5�K��`SKCFMAP  V�Wp�RM��M�����ONR�EL  lu�ơ�`��EXCFE�NB��
ģ���F�NC�
�JOGO/VLIM��dsa�.��KEY��d��r�_PAN����b���gpT�d���SFSPDTYP8����SIGE �����T1MOTV�����_CE_GRP� 1�V�ƣ\M�	�_a�M�Oό�mt vϷ�n����Ϥ���� !�G���k�"�dߡ�X� ���߾��߲��1�� U��_��r��f������	�J���QZ_�EDIT�����T�COM_CFG 1����h�z���� 
I�_ARC_���vD�T_MN�_MODE���@�_SPL��&�U?AP_CPL��'��NOCHECK {?�� �� FXj|��� ����0B�T�NO_WAI�T_L��>�)�NU�M_RSPACE๯ �����$ODRDSP����#��OFFSET_C�AR4�&DIS�/#S_A��AR�K��?�OPEN_FILE2 ����?���PTION_I�Ou�ɱ� M_PRoG %�%$�%��/�'f#WOR ��9�ԡ  ���6M�=�M�Ӡ�� �M� 0� 1	� �K� 1M�s���RG_DSBOL  wơ����?�ORIENTkTO��M�C�Ȱ�šA "U��IM�_D�'â 2�V~�LCT ���9�4�M�d9�3_�PEX��5/0DRA-T�� d#�0D �UP ��>p�>���O�O�O�O�I�$PARAM22������$�3\"@�_ 0_B_T_f_x_�_�_�_ �_�_�_�_oo,o>o Poboto�oM�2_�o �o�o�o�o!3EW'��o���� �����#�5�G� Y�k�}�������ŏ׏ �����1�C�U�g� y���������ӟ��� 	��-�?�Q�c�u��� ������ϯ���� )�;�M�_�q�����h<p��Ͽ���π)�;�M�_�qσϾ� ���\  ��  ��  ���  A�  Bl��4�B��C���H��&0������B���z��ͳ0�1�hP E;� E@ D�����D����������  ���/�E��,�N�c�gP�E(�E�_�^�Z�m���J��Fҋѓ�/|עޯ� ��~�G�o�o���E�b�D�����c�cќPЛ��M�PU�C��M�W�K�k��o�C� W�k�k�K�C��[��
o�m �NP�W�o�K� ����o�W���n���V�xԿ�+�I�C�U�0����І��ȍ��� ��k����k� Ћ�4K��ڌ�� ��������`����Fp EG�6#��F����c�g��@��������h	�����D��� %	GU��?��W%���p�O0���Ap����������./*$'� �$B��2.�� � |/�,��	�`��/�/�/�!:�o�1??%?7?@B�0N2��b&?��Z�����0D�� �� �k@�� �� �� J� f8����?��?�?�?� OODO�l�D�@OU��@�!�,!���T�"l�6 �"_�� @�?��>�A��?� �A��C�H����N;��	l�B	 � �@� �,�^t0���@��� � s � � �Rw H���9H�H����H`�H^_yH�R*L�OP�g_qTw CFPB�0BG�C4�T�@�_YS��9�� ��k�ô��G��Q�_�_�_�8C�B<��=�RQ��)�_@ ��1oRP�Jc��9�?2\S�o_�aЗf7O��oXU	'� �� �bI� ��  �!RZ=�����o	{[R@�%ppn�AI�+�B�b<boTZNS0�  #'�v�Q�PB���R��P�R�_�� �� � }��QCW�/� &=^;?�TXB O�O5�-K06qw� �2O��.O�����Ϗ@�e5s0�`��.$� ,RR:�����FQy0Ib�?�ff0fU�g��� � ��Į�\Q8RPğҚ?�"��ASZ(RP �P 	�$�DQ�C�Dis����v!;�x5;���0;�i;��du;�t�<!C��7_t����D�C|�BK0?fff?6p�?&��XT@���A#ǡ@�o[ϥpi����w �E ��G&����D��[�F� �j�����ǿ����� �!�3�
�W�B�{����t���p�E�C	�X����,��%�� I�4�m�Xߑ�|ߎ��� ����]?�w���O�� ^�υ��ߩ������ ~������9�$�]�H�4��l��!A�� 
"��C{���w�r�>�t�?��Nl9pi��6s�Wa�C����` Ca�^K�(�( '�@�I��~��bC�@_;CLn�B�A�Q�>�V�È�����Y�\���
�YS��Q���hQ�@�G��B=�
?h���'T ��W����ɰ�B/�
=�������=cK�=�J�6XLI�H��Y
H}��A��1cL�j�LLPBh�H:��HK����	bL ��2J��H���H+UZBuc/O/:/%/^/ I/�/m/�/�/�/�/�/  ?�/$??H?3?l?W? i?�?�?�?�?�?�?O �?ODO/OhOSO�OwO �O�O�O�O�O
_�O._ _R_=_v_a_�_�_�_ �_�_�_�_oo<o'o 9oro]o�o�o�o�o�o��o�o�o8#yG�y�>D C�a��>l Ĉ����OCVF���z<���K�	�� 
E.�1��|�z(�_�h~��7�����'u�N��۟�����3lC�8ˏݏ낢���	���t�.3��}�#�5�k���q'�3�JJO�O���@}�����ןŜ Po�	P	�$�%�2���>�0h�S���w�������ү���{���  fU�ͯV�A�z� e���E��ѿ����㻃����;�)�K�)�ZK�]�  ( 5��y�s��ϯ������	���  2 �E�x���E�L�n3���q��B���,��pC�� ����@�}ߏߡ߳����������$�6�H�Z���?�q���������������
 a���������� �0�B�T�f�x�����خ��������V{�H��$PARA�M_MENU ?�O�� � DEF�PULSF�	W�AITTMOUT�RCV% �SHELL_W�RK.$CUR_oSTYLF�Q�OPTg�gPTB�|vCLR_DECSN ������ �!3\Wi�{�������S�SREL_ID � K�g���US�E_PROG �%��%�M/�CC�R) "g���`'_H�OST !��!e$�/Z*T�l/�#ą/�!�#�/Y+_TGIME'&u%��?GDEBUG ����GINP_FLcMS�%>S8TRa?�R7PGA0 B<��;CH`?Q8TY+PE������ O@O;OMO_O�O�O�O �O�O�O�O�O__%_ 7_`_[_m__�_�_�_ �_�_�_�_o8o3oEo�Wo�o{o�o�o�oT5W�ORD ?	��
? 	RS�0c�/PNS�u`rsJO�d�TE� COL�u�hOZ�7L)  P���p��u%d71TRACECTL 1�O��  {� "�%�"��|�v_DT Q�O��p��pD � W� z��p�q���ߍ��p߫ ��	�
�������� ��*����dВ���s��s	�����������X��!�"��#�$�%�&��'�(�)�*�+�q���r�q �q|��r���r<����r�������#��*C��K��S��;�,�U�3��;��C��K�U�S��[��c��k�U�s��{�탄틄U�C��K��s��{��䃄����� V*�W�X�Y�r���[�\�]�^��_�`�a�b��c�i�j�kP�t�����C��K���C����T��;�Ҫc����S��C��K��3�<��c�
�� .�@�R�d�v������� ��Џ����*�� <�N�`�r��������� ̟ޟ���&�8�J��\�n���� de�e*e�fe�ge�h��ǯ �q�5�G�Y�k�}�� ������������� 1�C�U�g�y������� ��������	-? Qcu����� ��);M_ q������� //%/7/I/[/m// �/�/�/�/�/�/�/? !?3?E?W?i?{?�?�? �?�?�?�?�?OO/O AOSO]E1�O�O�O�O �O�O�O�O_!_3_E_ W_i_{_�_�_�_�_�_ �_�_oo/oAoSoeo wo�o�o�o�o�o�o�o +=Oas� �������� '�9�K�]�o������� ��ɏۏ����#�5� G�Y�k�}�������ş ן�����1�C�U� g�y�����sO��ӯ� ��	��-�?�Q�c�u� ��������Ͽ��� �)�;�M�_�qσϕ� �Ϲ���������%� 7�I�[�m�ߑߣߵ� ���������!�3�E� W�i�{�������� ������/�A�S�e� w��������������� +=Oas���������$�PGTRACEL�EN  �  ��� ���_UP �/���,4�-�_CFG7 �,�-�YYs~|~  �~�ADEFSPD ��L���� INDTRL ��Ll8��PE_CONFIH}�,�,rY~� LIDE��L	0)LLB �1�' ���B�  sB4#~ u%�*�/�%� <<7 �?��+�/ �/�/�/)??1?_?E? w?�?{?�?�?�?�?�?O0J�"GO>OPO}O��/vO�O�O�O�O/)G�RP 1�d,��y"�  ������A�PH���@3R��A~ D�	� Ap�	@�� d�$VYfY'!' ��P �O�/O!�^´�S�_�[B�P�Q�_�_�_�_�_o/b��BC5;oto�npo <�o�a�o�o �o�o�o�o	�o-@f)v��APz�s�� 
����(� �L�7�p�[������ �����ُ���6��J�)� )
V7.10beta1�� @�{@�A&�H#Qjo�CC� B���oD1� ��C�@����� D���A@ #QB  HP#Q3C
���� AA#C��˕/b�-P~! ��)Eן-PHS3b~!�9�ÑG�B���B
ff@�33cB� `�AB�]�����@�����ӷ�Ӹ���{��,�o(� .f������ٯï�n�0���!�A%"m`��]� ,"T�f�!p�,Q��lGR8� B�B������BHٳ7�� �� õ�'�7�X� ,� ^7�������{�<\�;IS�;{�Io��YC��fW��s3B�33Cϑ���*o�kGQA�������g~��ą������HP���߲���A4$KNOW_M�  �T4$SV� �d)�%�r߄ߖ�����@�߷���Y^]3#MS��H���	k�����\���*lI��$�@�p�������@4!MR
S�&�T+j<���X���s3e���MOADBANFWD(��2#STQ1 1��,a�4TO�OL f�.c@P����
����B��G�s3Ga?p3GE��}��2�������	�ZERO������%(i ��4�+=na s���� ��@6'l��^�2i��2�4Q  �<�ze�3�����^�4��//^�5 6/H/Z/l/^�6�/�/�/�/^�7�/�/ ??�^�8/?A?S?e?^�M�AI�_T�3�O�VLD  �;�U��O`�PARNUM  l�C~�UOn[�SCH�9 �5�
kG4AyIW�EUP�D4OE>��U�N^�_CMP_��0m�X��'U��DER_C;HK�E��U�>�V�O
[RS��L��'_MOI�lX_Y_��_RES_Gh���;
ɒ�_$��_�_o ooIo<omo`o�o�o �o�o�o�o�<�S��\�_�o�U�5: �S5 Uty�S� � ���S� ����S .0�1�6��S�0Q�p�<u��RV 1�o�R�2��[�ToRT?HR_INR���1��U�d�MASS6� Z�MN��#��MON_QUEUE �l�U�}P8�� �N�@U6QN83�\�r�ENDx��_җ�EXE��q��@�BE�����Av�OP�TIO�˞PROGRAM %V��%u���ZOt�TA�SK_I�4��]�O?CFG �V�O�J�}�DATA��ֆ�װ
� &� 2 8�9��C���C���E�EB�B�B�������4��� w��0 Qw�Z�P�g�U�)a�p�
m�
�^� ��V�`���`�L��@�� Ÿ�����������|�/INFO��ʭJ��MOR�d�vψϚϬ� ����������*�<� N�`�r߄ߖߨߺߵ�5I"��ʬ �i|�6r@K_��ӆ�B���ENB�0��-�h��7���G��2�� X,		@Qo=���¿���$w�@Q���ӄ���_EDIT ������y�WERF�L׃[�RGAD�J ���A�  ^�?}Pj��B�v����:E��?ޠBz�ڠ <���KI%DIAG�����J!I����2٬��4�	Hm�l�F�ւBp`�UU�@ޡ:*N /P **:YI[�{�D*P`����8b �?��:Eω�B*8`��: ����܁*���A��;�GY n�������r�/`/ /�/<A�!.'A��,- �/z/�/?�/?�/�/ �/r??n?X?R?d?�? �?�?�?�?�?JO�?FO 0O*O<O�O`O�O�O�O �O"_�O____�_ 8_�_t_n_�_�_�_�_ �_�_�_fooboLoFo Xo�o|o�o�o�o�o> �o:$0�T� ���������2(	����8�ʏ���t$ ���������=�O�|�PREOF ڌ�8���ҔRIORITY����F�MPDSaP �4�⪗UTh�|*A�ODUCTe����R���OG��_TG1�j�����HIBIT_DO�2�5�TOENT �1��� (!?AF_INEԐ��>��!tc1 ��>��!ud���?!icmѯ��XY������8�)� fF�X�8��@���d�p����� ѿ��ʿ��+��O�@a�Hυ�lϩϻ�*���ތ��%i����^��?5�!Df!/p��b�5������|�:�,  肐��ѫ߽�����8��R�ZR�!�3�E�W�5����ENHANCOE �����A���dQ߷��  ʄ�k��s����F�PORT_NUMՓ�8���F�_C_ARTRE� +�>�SKSTAԗT�oSLGS���+�����Unothing����� ��������	�c�TEMP ����,a���_a_seiban&��"� ������1 U@R�v�� ����/-//Q/ </u/`/�/�/�/�/�/ �/�/??;?&?_?J? o?�?�?�?�?�?�?O �?%OO"O[OFOOjO �O�O�O�O�O�O�O!_ _E_0_i_T_�_.c�VERSI������P disa�ble��]SAV�E ���	2670H722�X	�_$o!��&o8o㯆\o 	�hޒc��k�o��e�o�o%�3z�l[of���W_�#� 1�+�`�pƅ7,���*�^d�URGEv�B)�M��WF�pI�ה����W������WR�UP_DELAY� �3��WR_?HOT %������'�R_NORMALu� ���ڏ��SEMI��ߏ�b�_QSKIP�s����sx�_c��_������ n���ҟ��ʟ ��$� �H�6�X�~�����h� Ư������ԯ�D� 2�h�z���R������� ���
�п.��R�d� v�<φϬϚ���������U�$RBTIF��[��CVTMO�UL�:���D�CR�s�A� {�z�CK����E�|A�PV�D8�@Z�'�n��R��Ţ�=1�¥�繟x���߳�;�x5;���0;�i;��du;�t�<!��������#�4� 4�Z�l�~��� ����������� �-��RDIO_TYP�E  �}�*�E�DPROT_CF/G �A�c�}t�BH�Ev�;�2��� ��B� ���������' K6��|��� �����B0 ft���^�� ��/�//,/b/ ��/��/D/�/�/�/ ?�/(??L?n/s?�/ D?�?@?�?�?�?�?�? $OOHOj?oO�?PO*O �O�O�O�O�O_�O2_ TOY_k_*_�_&_�_�_ �_�_�_
o�_.oP_Uo t_6o�ovo�o�o�o�o �o�o:o`oQ�x�?INT 2�x���=�BG;� ��{�������f�0  ��{�
)�+�=� s�a���}���͏��� ߏ����K�9�o�]� ������ɟ���۟� #�	�G�5�k�Y����� ��ů���ׯ�����C�1�g��EFPO�S1 1�G� � xSAF�E10 pal �load
彳����q@
��z5��>���6X{5�ٰ?��6o<��5���5�}���20 la�ser mark軵s���q>8��8X@�H*�M�^��>[�?�8���������3'�eak� L��5��q=��o%���#���ٳ?�6Կ8?K��(`�v�Ԅϖ�4��R��  ��q�1k�0�j��]�@l�苾�R;�
�����������5�0 assemb�ly!�4��/���Z*����?
N>���?�<RP�f�tߚ�6��un��7�4�?I�Եs�����������70 �conveyorus��̲a�,�p>�T�b��100.�'ste��6�4ҵ���������
HO�ME/PERCHO rac2�5�$���ԿVwP?�2��5�ɑ�2�0,��0�F�T�� MAtpE�NANCE��8�8����)�Ѱ62'�а�,�٨����� ��?e	/�
�e�| �P�t��!3 ��{�:� ^���/�A/� e/ /�/�/6/H/�/�/ ~/?�/+?�/5?a?L? �? ?�?D?�?h?�?O �?�?�?KO�?oO
O�O .O�O�O�O�O�O_�O 5_�OY_k___R_�_ N_�_r_�_�_o1oo Uo�_yoo�o8o�o�o no�o�o�o?�oc �om���X�| ��)�;���"��� ���B�ˏf�Տ�� %���I��m������{  ��2 1헿 A�S������/�5�S� �w��t���H�ѯl� �������Ưد�s� ^���2���V�߿z�ܿ ϰ�9�Կ]������ .�@�z������Ϛ�#� ��G���D�}�ߡ�<� ��`��߄ߖߨ���C� .�g���&��J�� ���	���-���Q��� ���J�������j��� ����M��q �0�Tfx� �7�[�| �P�t��!/� ��/{/f/�/:/�/ ^/�/�/�/?�/A?�/ e? ?�?$?6?H?�?�? �?O�?+O�?OO�?LO �O O�ODO�OhO�O�O �O�O�OK_6_o_
_�_ ._�_R_�_�_�_o�_ 5o�_Yo�_ooRo�o �o�oro�o�o�o U�oy�8�����3 1�ğn� �8�#�\�b����� ?���ڏu�����"��� F����?�����ğ _�蟃����	�B�ݟ f����%���I�[�m� ����,�ǯP��t� �q���E�οi�򿍿 ϱ�ÿտ�p�[ϔ� /ϸ�S���w���߭� 6���Z���~��+�=� w������ߗ� ��D� ��A�z���9���]� �������@�+�d� ���#���G�����}� ��*��N���� G���g�� �J�n	�- �Qcu�/�4/ �X/�|//y/�/M/ �/q/�/�/?�/�/�/ ?x?c?�?7?�?[?�? ?�?O�?>O�?bO�? �O!O3OEOO�O�O_ �O(_�OL_�OI_�__��_A_�_e_�_��t4 1���_�_�_eo Po�o�_�oHo�olo�o �o+�oO�os  2l����� �9��6�o�
���.� ��R�ۏv�����ԏ5�  �Y��}����<��� ןr��������C�ޟ ��<�������\�� ��	����?�گc��� ��"���F�X�j���� �)�ĿM��q��n� ��B���f��ϊ�߮� �����m�Xߑ�,ߵ� P���t�����3��� W���{��(�:�t��� ��������A���>� w����6���Z���~� ������=(a���  �D��z� '�K��
D� ��d��/�/ G/�k//�/*/�/N/ `/r/�/?�/1?�/U? �/y??v?�?J?�?n?��?�?Ood5 1�o�?�?O�O}O�O �?�OuO�O�O�O4_�O X_�O|__�_;_M___ �_�_�_o�_Bo�_fo oco�o7o�o[o�oo �o�o�obM� !�E�i��� (��L��p���/� i�ʏ������6� я3�l����+���O� ؟s�����џ2��V� �z����9���ԯo� �������@�ۯ��� 9�������Y��}�� ���<�׿`������ ��C�U�gϡ����&� ��J���n�	�kߤ�?� ��c��߇��߽��� 	�j�U��)��M��� q������0���T��� x��%�7�q������� ����>��;t �3�W�{�� �:%^��� A��w /�$/�xH/.O@D6 1�KO �/A/�/�/�/�? �/+?�/(?a?�/�? ? �?D?�?h?z?�?�?'O OKO�?oO
O�O.O�O �OdO�O�O_�O5_�O �O�O._�_z_�_N_�_ r_�_�_�_1o�_Uo�_ yoo�o8oJo\o�o�o �o�o?�oc�o` �4�X�|�� ���_�J������ B�ˏf�ȏ���%��� I��m���,�f�ǟ ��럆����3�Ο0� i����(���L�կp� ����ί/��S��w� ���6���ѿl����� ϴ�=�ؿ���6ϗ� �ϻ�V���z�ߞ� � 9���]��ρ�ߥ�@� R�dߞ�����#��G� ��k��h��<���`� ����������g� R���&���J���n��� 	��-��Q��u[/m$7 1�x/"4 n��4�X �U�)�M�q �����T/?/x/ /�/7/�/[/�/�/�/ ?�/>?�/b?�/?!? [?�?�?�?{?O�?(O �?%O^O�?�OO�OAO �OeOwO�O�O$__H_ �Ol__�_+_�_�_a_ �_�_o�_2o�_�_�_ +o�owo�oKo�ooo�o �o�o.�oR�ov �5GY���� �<��`��]���1� ��U�ޏy�������� ��\�G������?�ȟ c�ş����"���F�� j���)�c�į��� �����0�˯-�f�� ��%���I�ҿm���� ˿,��P��t�Ϙ� 3ϕ���i��ύ�߱� :�������3ߔ�߸� S���w� ����6��߀Z���~����8 1�O�a��� �=�C�a���� ��� ��V���z���'�� ���� �l�@� d���#�G� k�*<N�� �/�1/�U/�R/ �/&/�/J/�/n/�/�/ �/�/�/Q?<?u??�? 4?�?X?�?�?�?O�? ;O�?_O�?OOXO�O �O�OxO_�O%_�O"_ [_�O__�_>_�_b_ t_�_�_!ooEo�_io o�o(o�o�o^o�o�o �o/�o�o�o(� t�H�l��� +��O��s����2� D�V����܏���9� ԏ]���Z���.���R� ۟v�����������Y� D�}����<�ů`�¯ �������C�ޯg�� �&�`�����忀�	� ��-�ȿ*�c�����"���F��ϵ���MAS�K 1�������!���XNO  �� �&�MOTE�  B���x�_CF/G �������A��*SYST�EM*v�V9.3�0162 ��9/�2/2021 �A �����R�EPOWER_T�    $�FLAG������START �� , 	�$DS�B_SIGNAL���$�UP_C�ND9�  �R�S232�� � �� $COMM�ENT $�DEVICEUS�E9�PEEH�$P�ARITY9�OP�BITS9�FLOWCONTRO8�?TIMEOUj�;��CU��M9�AUX�T��:�INTER�FACx�TATU���_RAP�C�H � t �$OLD_~�C_�SW ,�FRE�EFROMSIZ���ARGET_�DIR 	$�UPDT_MAP����TSK_EN�B�EXP?�$�!�o�FAUL"�EV��P�P������ !c�$U�SAGE�ENA�BL��	�IN_E�X��IO&�E��Y\��2�_ON�P��\����WRK�D���_TYP����IN�DX���������F�RIEND_GR�3�$UFRAM�_NUM&TOO�L0MYH��&L�ENGTH_VT�EIRSTX �#�SEF�g	UF�INV_�����$M�I��$W�AITING]
X�2l�G2��G1�������PRE9_+�NO_v�#��I_REQ�Cq�1����C3�n�>2A�GP_���� @ ��v�	�� ����1�  �E�d� �s�X� ��E_Me�CT��H_������Jq�G3�W������DEADLOC}K�DELAYE�aT�!$�$KO 2����1���1����2��2[+3��3��K)�!��i)�!`�������$V�ZnV�V3l J|�� � ��
4#M��h��.;"1PS��z��Z2�m���lACp9P#RDq8��#S� ;��4��o�Y� q0#��@  6!I2��q�� ��l � 
�q�S��	 �1R?���M�[RUNN��A)X��A  LT�^)BTHIC��	��IJ���FEREN|�1&EIF_CH���)AI��sC���0G1��8�D��IA�n n�F_JF�GPR3 ��0	�RV_DA�TA��
  �$�@E�� @� 	_$VALU�A�H�# _ ��A � 2
 �SC���	� �$I�TP_�B'1 " O9UQ1CSTOT DCS�DSPZVJOGL9I�� E_P ��)O:A=S� X1 ��=K:�_MIRvQ�T2� M��UAP�uE���PA�EQ�ЭQ9�vEQPG�VBRK�@�NC @It1 � b��bER$0ADxx�CS�PBSOCNV�x�NJeDUMMY{16�1$SV��DE_OP��SFSPD_OVR���0c�LD�b�SOmR�gTP@�LE�f�FZA�fsPOVvUS!F�j@�c�F�f:���S��h:9�LCH�DLY�WRECOQV�d,�sPWe Ms`�;uvPRO��Va�P_\@M� @��S�@�NVER��,�OFeS� C PWD�a�7t�aVa���Up`TR�8��Q�E_FD}O�VMB_CMQ1�pBfPBL%2�R�r%1�4V���,�[0;S2�bG�w�XAM�S�p0���^r9�_M�p���M:P��jqT$CA�iPe�Dbp�HB�K0�?���IO��2��I��U0PA�������Ą��D���jsDVC_DB���@�+� ��Gr:�����^��y3�dpATIO�������aU��hPh���ABP����Hs�����sP_��?�S�UBCPU*�PS ����s�1��ȗ�#��
��1$HW_ACK ��"#��1#A�~�0�$UNIT'd�!��ATTRIxB�.��PCYCL���NECAZ��SFLTR_2_FI�D0?�`�1��LP�[k@�j@_SCT�F_��F_$���6�FS80��r�CHA��p��r���RSDhp`,�7aJ�+ᬀ_T��PROF��s��EM�P��vPcTۢ�!c ۢ�a�DI��~A�RAILAC�eM,PLO:`Lbd�5&W0d�_1d�^�P�R��S4��̱C��k�	]sFUNC�2l2RINS3�-��v�촭�RA��1 �p��;�~��WAR�Cq�BL.+�F�aA?�;�B�;�DA%`0���F�?�LD!�x`����!A�V1��TaI^2��>Q�0$t�gRIA�:�AF��PH���Vp��h "��|�MOI%��vD�F_R �c-��LM��FAe HRDY.��ORG��H�3�-���G�MULSEPR B�ȗ�!n�J�j�J�b�g�kFAN_�ALMLV8���W{RN��HARD�� 0�d�L� �2�ѓ�d;Q�U_2p?�AU���R���TO_SBR�0�gP;������S�MPINF@p0�f��q�REG��cNV.��fDA= ��tFL���2$M x�kE��^������CMf@Ni@Y�NON�p�{`G�p�p�.Q �0��$.��$Z�*RQ�/P$ ��SEaG^0CSx`S�ARUPi�`e27&b�l��UwAXE]WROBZZ�REDZVWda_��<cSY$`��`��S��WRIe f����STRYU1�`�`E��@o�8jb�o�B m�%9��J�O�TO���@VpAR�Y C\��J�Q�QF�I�P�S$LINQK6�0A|�!_�m�ad3�0��X�YZ�Ү
��OFIFrp{��` 	BXP�Gqp�FI���1{bpd�rT_J�Q�B�b����4>
3�F�TBR�ҊCp�&�VDU�r`e3�1��TUR��X���jba�X��e�rFL� @py�`���!	3ic^�q 1�@KPMd���ȕ^2ȗ�s�ORQ>�gQ�x6 ���P�@8�_1�%ceQ���$OVE�!3BM ���A'��%-��%3��& ���({��'��$�E� ����4A�!�P0��A �%�!�'P5-�P5�#gQSER�Q�	��E��H�@���4A<1���9�h������AX Gs�B��5��}�5i� �9���9i`�:���:� ��:v��:. �:L �:1 � �6s��9s� Is�I s� Is�0Is�@Is�PI s�`Is�pI�A�I_�6���5DEBU�$����a�AQ�r�AB������a�#Vz�� 
\R�h1�U⑐W ��Wia�W���W�!�W v�W.�WL�ď��\$2LABr%���GROs�r��c�B_G�u6
B� 8�9fmas%ie&�ufAND/ ���4d���1&�g c��� �h0x��hf�� NT��;s�`VELM�"4q��
xQzNA���C��c�v�$.���SERVE�`�B� $��;q!~pPO����p�V �qOmr��A�v�$�rTRQ��
�s��p�w��2��v����_  ql�0�є�ERR>�i�Ie�p"4�TO	Q"40L���4��&��9�G�u%���� ��sRE��  a,|q�u�p%2RAh�? 2 d����sTc��p "�$� L�)��27�q�OCx��p  }�COUNT�_�lpFZN_CFG�q 4����l��T���3�5S1q3� �MIN�>� ��P5�T�/343�!�\�FA��-5��`�X����\�<�g2��ҁtB���P��_��SHEL����� 5JB_B;AS��RSR��հE��S����1O���2�3�4�5*�6�7�8O���RO-pU�� � NL�-�AB�s��A�CKmVIN��T_���U�~�ࡡ�_P�U�����OU�sP�8���ΓP�*� �6T�PFWD_KAR�����RE�t]�P8x ���QUE��0 � �����I��pS�Γ� ��p��SE�M����=�AX�S�TY��SO��D�I����.c\��7'�_�TM��MANRQ�� END�$�KEYSWITCaH���ϱe�HE��BEATMG�PE�}�LE��U`E�U��F���SԴDO/_HOM��O�Ѥ�EF� PR ��� ��C_�Oi��h�OOV_Md��EGOCM�l��wPv͕HKA� D�$��.�U�rZ�M[�.��� �FORC��WcARYҿrϓOMd�  @KT7%�UP|�1a���c�E3a�4ha`���O$��LG�q���UNLiOڠ�t��ED��  �SQ`HD�DN�q �pB�LOB  ���SNP
�S�� �0��ADD.�0��$SIZ��$V�As`Q�MULTI�P����f�AG�? � $���H����S.c�C��`�FRIF钳�S�D�Vٗ�P�NF�ODBU���`n���X�v���IA5�Ac��8&Zx"6��B�� � 
�0�TE��_r.SGL�T��&�5�:c����STMT�N�PS�EG��BW� �S�HOWV��BANb�TP� ZwL(�h_s�̐V�0_G@�;  . $PCB`����3�1FBC�P��S�Pl�A������VD���?�!� ��qA00Kuj�$@t�$~�$��$5"	U6"	7"	8"	9"	A"	B"	U�$a%�=p$F"�@�.	1P;	���U	1b	1o	U1|	1�	1�	1�	U1�	1�	1�	1�	U1�	2!	2.	2;	U2H	2U	2b	2o	U2|	2�	2�	2�	U2�	2�	2�	2�	U2�	3!	3.	3;	U3H	3U	3b	3o	�Xp�(�	3�	3�	3��	3�	3�	3�	3��	4!	4.	4;	4�H	4U	4b	4o	4�|	4�	4�	4�	4��	4�	4�	4�	4��	5!	5.	5;	5�H	5U	5b	5o	5�|	5�	5�	5�	5��	5�	5�	5�	5��	6!	6.	6;	6�H	6U	6b	6o	6�|	6�	6�	6�	6��	6�	6�	6�	6��	7!	7.	7;	7�H	75Y7BY7OY7�\Y7iY7vY7�	7��	7�	7�	7�	7��Ip��PC�U�rQ"�ҡ`�
��V���uq# x $T�ORM����Ђ��pRX�p���dQ_̀RrpP(��q�D�S�mCo�u v_Uy�+q*��YSLM�vp$ � 
��������y���0r�Wt��VALU��Ơ��a�xFHqIgD_L�uHI�z�I5�$FILE_X��t��$��ADu{SA��% h�`~�E_BLCKG���7�%�D_CPU 5��5������t7��Y��R & � PW΀����6��LA\�Sǀ��\����RUN��G�� �����Ņず�あ��H砱����T�2�_LIG�' w ��G_O��}!�P_EDIg�f�`T2u�%�(-��ٙ�0�R���O�T�BC2) �������.�%�FT8������TDC��<�´�M�஖đ��THD��g�ڔ�c�R��<Mp�ERVE���������y���ݐ *X -$3�LEN��@���3�ʠcRAC���GpW_q�b�13��t2z�MO$-���S�๠IϠr`�q���d3���DEǥ���LACE���cCqC��rW�_MA��pƦ �֧ �TCV�(�֧T��)�H�>��� ţ��l�֣��J���`��M��M�J߷ ť)��֥?�2��w� ˱ģMpJK޶V�KG��������Jخ����JJ��JJ�AAL��*���*��$��(�5�[�N1�O�[���tL��_dJ����/�CF���+ `�`GROUP�p8����N��CH�~��REQUIR󒎱�EBU_�/���$TǠ2*��0���8y����, \-p_�oAPPR��CLr�
$6�N)�CLODk�9�SЕN�ť
y�.3�- ��M�8Z��҉�_MG��ЁC ��ؒ����B{RK��NOLD��}�RTMO$�������J$���P,��������H��Q��6�7�*��/��.� ��Z�G��y�����PATH �����_���y���9-q��SCAc���l*Ғ�IN2�UC�������C��UM��Y|�����q������3��PAYL�OA��J2L�`R'_AN��^�L��h��d�X�t��R_F2�LSHR���LO�i�@�������ACRL_%�������P�r��H�pr$H���FLEX,�X:y�J}�/ PҎ����������J2�0 :?�Q�֠���T�S�֠]�o���F1�������Ưد�KE����*� <�N�`�r���"(?$�� ��޴/Q(����ɿ�кT�' !X(q��ܵ �v��%���� )�-�6�$�H�Q�c�u�t��,�J��1 ���`�Ϲ���ؐ�`AT4����EL��C�ȵJ��0��JE��C3TR��/TN�aF���HAND_VB�r,�pm�2 $�� F2��Ҕ�sS�W,+�w�3� $$M�����`�ѳH@���L��E��FA�p U��־q�I��A�܁p
��A��A��	P��N����D��D��P��G���YST�קQ�٧QN��DYĀ'Н��D Uv�4��������W� ޷v$� � ��P!�*�3�<�E�N�W�`�r�J�~�4 �@��� �\�e[ѱaASYIM��p����3q�����_�����
� ���dzH�&�8�J�\�Jc��u��s�y��A_VI]C�x[��pV_UND��p�s3��Jߵ�>e���� ��!�E��������������#%R 7�T��HRm�b��5sBƁ? 9�DI$����O�Ѱ�Ɓ�ç6 )0RI�aA ����5 s �8u��K�7Ȁ 7 �[ �AME�m0h;���"qTـPTxp �0��c�����> Zp�h���w�Typ�� �$DUMMY1�3�$PS_2RMF�   �ྖ��7FLA��YP�#ؒ�k�$GLB_T`�@ۅ�c�GO�p3A?�8 X���m��ST����SBR���M21_V��T�$SV_ER��O��09�Q�CL��9�A��O�GL�pE�W��9 4��m�+$Y2Z2W��԰���CA<���aB~�U.��: � N��~p�$GIC@}$>�� 9G|������; L��צLr}�$FLrEߦNEA�R�N9F&��T�ANC9�JOG�� 
� <� $JOINT�!��q��~�MSET��= E ԧE�6�0S�2�_��0��>� � ;@U�?���L?OCK_FO��A��BGLV6CGL�иTEST_XM�,Џ�EMPb���8�����$U� ��F� 2:�����;�h�@���9;�CE��|�;� $KAR�}M�TPDRA��X�O�VEC� i�S�kIU�<�HE°OTOOL���V�;REp�IS3z��96<�/ACHu���E=��O��k���3���SI�  �@$RAIL_B�OXE�!^�RO�BO�?�^�HOWWAR
ѻ���ROLMƒ0Ֆ1���A��1��#o�O_F��0!^�HTML	5ځ���5�@�2��-GC�CHp�?[���Rs�O�@[�� d��hЉ~�OUw�A 	t^��9"qB�1�����PO��@PIP�N� ������A���� CORDEaD�����#�XT	�ڡ)�P�0O"� �B D �OB>QC��i�X᧓�X�LpASYSX�A�DRAc�TCH��@ C ,� E�N˂HAǱ_פ���1���VWVA~>�D � ^����ۅPREV_R�TKa$EDIT�
�VSHWR�1P%�)�����pDM��@�1$HECAD]q��Z�mq��KE����CPSP]Dq�JMPu�Lڅ2�R���E`�=���I��SBCW@N�E��AMGTICK��sqM�1�1��H=N�F @b���5y�_GP��I gSTY����LO��k����@G��
��G��%$��פ=:%�S0!$�� �R�ޕ�ݖP�`S�QUR��ߒ�qTEsRCg�G��TS�4H ޠ1��7� �7R!��@Oh�[�=�IZ��סܕ��P�R;�Ǒ&����PU��q6_DO+���XuSs�KچAXIUT��UR�0�B �����A�0_����ET�Pɲq��e�T F�gU A�Q�a���9��)@���L� RjDIl � �I�"�J%�F#)�B %�G#�I#
YW%,W W%<WW%LVi%�-yYi%H�,�b�)C�/�-C�-�EWi{t��SSC��� J h^�D1S 񁭐SP��5AT:P�B7����~��ADDRES��=B�SHIF����_2CH@�I\��1�TU�I�A� K[�CUST�O��AV��I �L���ݸ�1�`
��
���V��F@�M \�����T %L�� bBCxS��4J��W�bA��TXSCREE�Z�NҀpTIN!At�堵Dפ���2�`O T��T� ��S�0�Vc��c�D�RRO`@���k���A{?UE��P ���`��̐Su���RSM��YUD�� چlQƀS_���V�c|Q�Y�W�c�C��hR�DO 2OJR�dQ��d��V&GMTX�L�2�r@� �h�� B�BL_��W��O@RS �T ,bO��8b�LE�2Cc��2BdRwIGHLcBRDf���1CKGR��teT�E�sgpaWIDTH���6�z��ؑ��L7�UIc�EY~�?�S d��s�/�8��="BACK6ƒ4�ej�F�FO2��g�LABA!?(F�I<����$UR�'p� 	�aL�H"Q 'T 8��@�_Y��2JrM�R������ȶ���07qO�1O@U��$q�m`UX`�sRɲ;��LUM�sz�0ER�V��@�`P*��dVD��GE+r��LK�b�LP�u�E� H1)�g��h1�����5�6�7�8 �r�!*�vD�������S� U�aU{SR��W <��bL�Uۢ
CۢFO�0.ۢPRI�m����TRIP��m��UNDO��XҠy �["�Z�p8���  YEr��.%G a TT�61L�1@�OS��U�R�(R,����QZ�������|�JQ�U�q�Q[������S�r,�OF�F갇�\z0��OD��Z^����[^�GU��P��8�31�B��aSUB �TE_EXE��V��,�WO,! ]2̐L�nWA��w����0V_DqB����3rSRT~���^��?�`�OR���ޥRAU
 ߤT�����ġ_��_ 9| ��OWN/���$SRC3P��w �D�J�"MPFI8/N1�ESP2� �@���s���w��+��#��Q` `ΐ������ COPב	$�1�_e��ر��ߵ��CT�c�������®���.�A a~�BSHADOWw���.�_UNSCApw�.ìd;�DGD���p�EGACҳG_��VC9 Cœbǔ ��$��ER�@�̙���yC�Л�DRIV�_V ����/��D��MY_UBY ����[|��4Q� �@bG�)��8�P_D��/J�L<BM?a�$��DEY��EXX��@S�MU��X?a��ԁPUS���_�R�A�ـ�04R�G>� PACIN�� RGT�������Ң��ҴSرRE_r�1|���������c �0ʰG��P�B"�t���Rl���d�`�p!Qd�ah�	ײSRE�ӛSW��_A��G�$��$O���1A�0��"EUG a�������HKLe�p��� !��P��EA����焠Lp��I�MR�CV�Qf ��pO*X MLpC�C	&����&�REFgH�/� ���p�mเ+�~�@<�~�M���/���_G������� S����������� ���Tg ��r��c�3Ł��� OU�0����� b8�712c`�P�@x@%`d�3�71j]P�0UL� �e��CO`Pאf��} NT���¾ yq����� L4���D��yq����V�IA��h �6`HyD�0�`$JO���b�$Z_USPL�9QZ^ WYp+�Rqb_LIfQ$EP}b�M�I +�A�1�v�0���OT�i 5�3PA��a �3CACHV�LOr������h�a�i�C�MI�3�F�"%To !&$�HOLp=��COMM��hROV`W'9��b�^��q=o�VPx�|�"_SIZV��$Z�Ъ(Y�'���c�MP�*FAIYG����AD�)زMcRE<2�'GPnP�v�^��ASYNB{UF�VRTDQ5�]4�!�cOL�0D_tݓy5W��PC_���Uo��Q��A5EC;CU�VEM���<�2 'VIRC�!q5�Y3gR]1_DELA`�^�3� �%�AGm9R��XYZ�P�S�сWS�1Hp�0D�a�0T��p�IMAp6�2�`�%GRABBy�Y\�ӟ�LER��Cr �F_DLЪpv5 �P�F��Enr����Tuj���bLAS�`\V�_GE�kWR^��2s3UTg^��������I9T��6���BGH`Vq��PK����6�9GIPN�p��k��B�,1�Pl���S!0�N�TC'�VLs��m)�� �qs����!�`Iw�C3@e��X4��Xf����(�1e��n���ZJ$�rt�����D݁��'ۀTb D	�o -$��IT��n��Q8�~���VSFͰ ��p  ����MU�RV��`M�9q�,�ADJ�`��v)ZD�fr DBh�zALc0�pyP�ERI�B$MS7G_Qq3$�!�%�@���	�s��gI�x���k �XVR��t�BD�T_OVR~�R �ZABC˥!u4�rJ#g�
�Aq�ACTVS� �v $�u�/rCgTIV��k!IO!Ҙ	�f&S�ITy���D�Vx�
���A�4�!V�D�PSde�� 3e�k!e ?�k!L�STS�k!q ��_�S���QqDCwSCH!�w L֡ ���u o�`�h� � GNAi#x���k!���_FUNc�k �Zd?��tx�Ru�$L���e��̒�ZMPCF˥y�b*����j�=���LNKT�
�)�)@̤z �$d!��B�CMCM��C�C˱~�T��P�q $J����D�!�������������;�B����U9X<AA�UXE��� <A�����������/���FTF���\��V��Z �{ A�k� Z� �Y�}D�@ | 8���R0U7�$HEgIGH�Ӟh?(� ċvf��@v�'} g� }��q$B� x��TŻ�SHIF�#��RV�F=pg���pC@��˱�~��� 5�W�S]��%Dm����CE��V2At�SP�HER�� ~ a,� ��ǯ٩ ���PL��N<p \��������ԲOWER �����SM_7DRY�% ��%��3�D��9��Y �N�UM�O� /Ϫ�� `���P��=�GSPD� �P�����_0����R�d ��I_AIR�PU;�  ��  �ϲ��0 ��T��p"ISOLC+  ��c�J�p'�����21��	�fu�?	��R��<0!T�P���b��3�;��t`d? ��`�H722  s�v���԰�0%�x԰S23�2� 1 ���� LTE� ?PENDAN��s����	�s���ϓ�Mainte�nance CoKns(��(�""��4�No Use �R��v�������������Nf"��������CH�Q 3����	A?!UD1:gRSMAV� �q��O�����P��1� 2�� 
PAL 1P���	��������2@Cz  D��� �N���a  E� D�T� < � ?��K�v$�{��1�4��Ăv#DJ����
�@ER MGARK��\���|0E0 C���e(!9� Dc� D�@BdZ/�`��/�/��L�G L/f���y�%$� �D �Dr` (!R�.B� F/h/^?�/�/�?�?�/�/�#R�/?�� ��D� ���67. ���F?h?^OO�?�?�O�?�?�"ASSE�MBLY�?O�!���#9�Z� �����G%  �;A �MOoOe_�O�O�_ؼ_�O�O
�UN �_m�\�*LQ,?/B�@:�S_ u_ko�_�o�o�o�_�^	CONV F� ��Oo�#��+Z&�9@C1'�` D�)/Uowom�o�o����o�o�dIMPQG�5��3~� F{�9@Xzp� ����Ǐ��� ����/�6��%7D~0�� �"Ed��  �*P EE/�u�Ϗ����̟@ۏ����?�
7��� %7û�J�N@ Z�|�r�������ɯ؟����2��  � �3���֧ g�����ٯ����ڿ��3�"�4�F�X� 
�|����������������41�C�U�g� y�+ߝ�����߲��)� �>�?�5R�d�v� �ߚ�L������9��� )�J�!�_�`�6s�� ����m����Z�@��JkB���7�� ��������� 25�{k�c��8 ������!S V/�6/�/�/�/�/�oG �At?r!
#0 ?  �C?U?g?y?�? �?�?�(�=��/�?�/-Or!dC@(?:?hO zO�O�O�O�O�O�?�? �>�J_.[K_>OPO�O �_�_�_�_�_�_�O�O __8_Joko^_p_�_ �o�o�o�o�o
 oop$o6oXoj `%$�ߩ@堣u�5�Ăt�DJ��H篱|L|�wz  ���z�%�g�y� ��M����ӏ������ �-����E����� ��m����󟽟ǟٟ�M��|
O��"��_MODE  x�"��S 	���GEz*/O���H�m�	h���G�CW�ORK_ADȬ���2�(�R  ���߰��ɰ_?INTVALȠ$����OPTIO�N � �I�V�_DATA_GR�P 2#x�D�`P~�j�z���y�{� �ϩ��������'�� 7�9�K߁�oߥߓ��� ��������#��G�5� k�Y��}������ �����1��U�C�e� ��y������������� 	Q?uc� ������ ;)_Moq�� ���/�%//5/�[/I//ϡ�$SA�F_DO_PUL�S��Р*q3�!� C?AN_TIMǡ�e�+��!R �"�"6��ՠYp!2'�A��q4��!�c ��1?C?U?g?y? �??�?�?�?�?�?	OV�jc@�22D$�!=Id2DMA��#I�p㾅O�O�O�B�aIuO W��D�_�t  Tް�O_�_0_=YT D��=_f_x_�_�_�_�_ �_�_�_oo,o>oPo�boto�o�!�sH��o�o�o�i  >;t;�o�dq��p��
�u��Dif�	1�j?� � �@�� ס	15�!t��� ������(�:� L�^�p���������ʏ ܏� ��$�6�H�Z� l�~�������Ɵ؟�@��� �2�D�����O m��������ǯٯ� ��L� E)�;�M�_�q� ��������˿б��0rWs%ua}�.�@� R�d�vψϚϬϾ��� ������*�<�N�`� r߄ߖߨߺ������� ��&�8�J�\�n�� ����������W�� "�4�F�X�j�|����� ���������0`BTfѿWq�op+�� � � � �mp�1����� �!3EWi{ �������/ ///A/S/e/w/�/�/ �/�/�/�/�/??+?`=?O?a?s?~7�o LS~?�?�?�?�?OO 'O9OKO]OoO�O�O�O�O�O�O�J�?�O_.)V���_�m�	123456�78brh!B?!�� rq�0p�_�_�_�_ �_�_�_oo%a�?Ho Zolo~o�o�o�o�o�o �o�o 2DVh y}7o������ ��,�>�P�b�t���p������{BH͏ ����+�=�O�a�s� ��������͟ߟ��<��{;�j!�K� ]�o���������ɯۯ ����#�5�G�Y�k��yD�u�������ӿ ���	��-�?�Q�c� uχϙϫϽπ���� ��)�;�M�_�q߃� �ߧ߹��������� ��7�I�[�m���� �����������!�3� E�W�i�(�������� ������/AS�ew������V����+=�YZCz  Aо�:   ��82�T}��J
��  	�J2�����R,?��P1�3 4 5 6/ [/m//�/�/�/�/�/ �/�/?!?3?E?W?i?P{?�?�?..P�2(�2 �?�?�?OO(O:OLO ^OpO�O�O�O�O�O�O@�O __$_6_=St�|<ZT PU~�  �j[��_=VgR��t C q�Y�_=X`���$SCR_GR�P 1"Y��"b�� � ��� w	 a�b(b!d	YQy>i�=W4gboPo�oM����bD�` D��@-.c�g�k+,�R-2000i�C/125L 5_67890��e~�RC2L p��c
V09.01 7pWhLR#� [va�fafca+#YQ�a%jZaly	]r������?��H�`�t�gvu E�y���6�7D����D���B�  �:ǟj���3aB� =�` �0A� �96GK�� S�JoY�>�(C�7�/D��]O�A`���oʏ�o�Sߌ�hR��Vvq߀  [_�Ǚ��B�  B�33B�=�D�<�M�3aAq_�  �aw�3a3@�u��� ?.����_�H=���b�3aF@ F�`ڒ�ُ ��*��:�`�K��� o���Si;��a��ӯ�� Я���S�&���J�5� n�Y���}���ȿ��� ׿���4�/-̰crodǉ�<i
�Ϻ��ß�@��.�4���Ã��`��=���1G234s!�x� P�Y�k�`�tՠ�Xc�P$��+!u҃ �߾����ڬ�������� �?G�Y�ߪϏ�z��@���o1Ԗ���qs��P�ECLVL  ΃��vr��+v���L_DEFAU�LT�����Y�HOTS�TR'�����MI�POWERF�xU3�\�WFDO(�� 3��QERVENT 1��T�� L!DUM�_EIP�����j�!AF_INEx'�����!FT����?!bWf��.�!RP?C_MAIN�nq�z��VIS��	��#!OPgCUA$J�o!TPbPU�f��d^�!
P�MON_PROX	Y���e�/�����f�S/!RD�M_SRVT/��gB/�/!R3Ի/��Yh�/�/!
� M/���i�/7?!RL�SYNpS?^78|&?�?!ROS���<�4r?�?!
C}E�MTCOM�?���k�?O!	�2C'ONSO��l
OgO�!�2WASRCdn/��mVO�O!�2'USB�O��n�O�O!STM��_��o�OK_Ro_b#<_�]���ICE_KL �?%�� (%SVCPRG1�_D�Z�U2�_�_�P3o o�P��4o�Q5Xo]o"�P6�o�o�P7�o�o��P(t�o�\9�o�k �T�/%�Q�_M�Q�_ u�Q"o��QJo��Q ro��Q�o��Q�o=� �Q�oe��Q���Q; ���Qcݏ�Q���Q �-��Q�U��Q�}� �Q+����QS�͟�Q{� ���Q���aˏ�_�R �P�_�Ph���o���կ �������A�,�e� w�b����������ο ���=�(�a�Lυ� pϩϔ���������� '��K�6�o�Z߁ߥ� ���ߴ��������5� G�2�k�V��z������������1��Z_�DEV ����MC:9� �CK�GRP 2���G��Pbx 	�� 
 ,��
���G� ��r��� ������������ Y@R�v�� ����1C*V�� HG��G��G�E;G���F3 y��'��/"/ 	/F/-/j/|/c/�/�/@�/�/�/�/Q[��� ��5r�/��U?<? 6;�?�/�?�?�?�?�? O�?�O�?_OFO�O�jO�O�OT�_'O�NG��O�O� @_�d_K_�_�_�_�_ �_�_�_�_o�_<o#o�5oro�N�G�MG��Dzo]f
Q^_�oZ_ �oZo,U<y `������	���-��o��D
G�6��G�f�i�o z?����ʏ��+� =�$�a�H�����~��� ��ߟ�X��֟C� *�g�y�`��������� ����ޯ��?�Q�8� u�\������Ͽ��� ��)��M�_�Fσ� jϧϹϠ�������� ��7��[߲�Pߑ�H� �ߜ߮��������3� E�,�i�P����������������&�d �VP]6t��	 ��>��V�1N���K����e7@�	�N{D�@�Y�����A�5��@*��Al2����|O_������E-3AyE�O@sž�tV�gB�uG_�?��>�����A�qF?��A���@�UU&�%�MOVESAFOE OS&���P;���?�?��O>��Kn>���>w�;#=P}ƾ
?����3C���Q,^����A�q{��w��@w�@.��3�� ��i����\�A���-A�XEBn��@3?�E���� �A�����V�AE/S>��3	��MARK�ER���RVP_�Z?��b�d?���J��)@B���	hZ��:<3@_<B���4>A� ?�	�?r�@�� 3>	������*���{�B�I�� �����Og3�ٳ���@y5@�~�A6����4^���ܫ��� DVP`G?���y?Q�:w��l?�!��5��L�A�3���b��ӐA���@}�@g�%2?��3������*�b���B�+o�����l^W��PmZ@����A��8?,4�-vy���v/�fy?�>W+�������Ύ���v�"?qk�P��4�W����s�Ԕ7?�p��@���4�3A��h�!���5�_�A![^C)�73�=�,@�����A,܂>;_��A�������S*APP_LA�SER���VPg�R?�=.~���7�*h�@����u�����3[�I�e��uAϢ�����rA7��@]�zE[8�B1����&0/B���AKjPC�"=�o��8�=CAL!:�C�.tA,�p�Y�y�S*ATTAUGHTPj!B?T;�m?�<2�����c��6Y�?������������W�zE���A�������AD�7@���?8�B1����'NvB��ALB�CP��>g�&t@ֿ��=y�����}50RO_D�EPARTO�H�_0r7F�m���x�d�>�����v���FZ�,B��N�Q#A�� �c��9A;3�@/�ƠO4�B4Z�]�.�B	��AReC������q�}��@�v���{A&��=%���K�_�Jl!�&S�ߙ=�^+4���W9@�%�@��k�3Kj�����A�^A���?�����3B��)��_�$A��B�&0�Q-B�Aͧ��(������@��s?��7�A[4�A��x�<60PALOLOADO�i�P�E���+�_K�n?l��>�������;���dy�� �HA����!���A]B?����nB�>�B���@��6�ǈ���v��B��*.�-E���z�qA�-O?19�,q��S/e"BLY� �`hptQVUm��?�A��\����+�V���NtA�p�A��^;3��o�h�0A�l�A��A�����"����.�׫���A��Uu;B��*�����<�ldS	����+&A(�H�^���Al8�@�ø�'?9?B�1@Un�1?�������U��Q-?��1^>�^�\�`1�������A�mC@�����F=@&��'n)��A��Q?��z@B�����'Y�Q�"��.0W����A$p���#o�?���Z%�d�UN�c��!VV�m�?�=�9���JA?�\�>g�)7�CN����6;�R�ĄA��rA�VrSArY�?���.��
�YP�A���
��!����B�,Oo�(�����A���^@%*@�7@̇�KzLe!�aET
��+���[�_�⼤��I<��@BD������^#�#-#�����A�a�@�2��1��}O�@��3���������B����	�H���j�/����$��_A���A���L �>��/ǟٟ�� �VVq��;i�@�jV@�Y�:A�����q��K�6�����D�A��F?"�At�?��p�.�3���I���d�B`����7��B�M��3�UB`��E�Aj��A1��y�,)R@�ó�Ke"����WV�V{<?�@\cO�?��/:�>��@5,������J���`�����'A��v�?�"�@���@>��'n��(��I?����BY ���-(�B��:���J@d@�c��@�b�@�7@ᾠ]|�a�h�AVV덏?�:P:&�{:%>�<:޼R����.���>���8A� ���bo���ߔA�3���;���F���CTo�i�T���d3�����Y��AI�.��V���C�i�-O�4�<�G{���7F�i>Y��]��"[�,N����,m���o�N$��8�A�խu?�x����pA<����a�?�<�!CU���`�a���>R*?���m���UA&��/�bi�1�*��V��^_LEAKTES�_��{�����_�;Dp������m�:o��AE�q/���lA�NA?h@��ΉcAA����������F�����c�iU������&����h�ATc���� <�m�@�@�&���JԎN?�;���m<��Q��c���Ϙ��+<U�!�N������A���?����tT�R\o��<�A�g����7�C@!7�?��O�>�r�X��@�@�^<1�?����_�_ܶ��PV�����_>�^C��3�F���� ��>9`3Q���g[A�^��?�����y��R�ZC�=��A�`���5�C@���x���>�اNI|�@�<�~������%��?DÅ�������������:�.�}���I>@���.@��)�D�N�4P���0�A��x�����>G@LP�o����m��OG.CK�q��Z�������@4q�
A!�ܾ���U��J>��b%�����a���r���>��_��_��>@��>�:�˾�ja�~��A�`@<��K;￥:��]�3��A�q3��o��B��������i�^�|�����A�>��A)��i��	��?F)/�T9V�ɫ��B����b�F�B���@�6y�@�J˾ ���˞A���A�ڼ�M�e���&:�"��d�)����}u�B��v�4�B���G����4A�qFA���0@s)��1�?1@W��ɿ�����]Y���:T@^�<�Bz�N� ���vAӳ9?��@<���w�'n�� �_0�A��_��0w0�W��d�8����A�H���Q��-ῐ�H�?�3jVX�k3���
}�9�-`?��AO����X�e���^i�,���A}����`�Alk'@�����]C�-�U���A|v���E���3?�CFG�'˾܁��%A��V@ ��A>ϭ�>x�� �CO?NVEYOR'/�H�	Vn|�/�����G���*����p�����?!>>�~3J����}�Aק?�@�P��<P��~MF��^	\���#�B�������&n�?^%%�;�}�@��@�Ś���1��:hc����߂_ Vn���[����?I�����@@zW�9���������~L�f����A��?����>�ք�Y�������������B����!�1_��as����q�)3Y��A4��7�a��l_Qo�V�&'��ň�?��$��;PJ@��r@	�>�~^�˾���L���sA��??K�h?���@Kj��� 0CA�#O����L�^-�A�/Ch��{���P�X%�A���@�(IA����9@o%,s�;k`Rֺ(0?KX�����?۰�?S`ۿ�R�G˾�<B����A��s��@�a�<�o#�A��ٗ�����T���A�=�Ce�η��ؗj�{�$PAH@���A0*H?�M��8w�/���&��<r�t�����<k$��s��} ^#A���m@�`A����G�q�C�A���*���n��O��A�ڃC�dY���G�:���^	A���@ئ�A+�3�8/͏5n����Lq�A>�x�A�:E���H���A`;�d�7�����A�e���*�A&S�@��rS^�L����v�'��N9A���C�Y6���HQ\x�A�[`A�A@�=�������n�ܛVʭr�A ��A!��>���>�[h^9������A�KM�?��:�R�����o����@��s��uo�CDXo��Ϸ��CB�˾L_���Q�A�����ށ��<-*���]�����z� �CVn�#�6���:T	��P��A�Y@hߖ�,����^[�C��z!_�����3�EN�@?�����$;��.[�](�C>���������˔˾��P��BIAS5�?��=��h�ڿYcyɷ?�?N� T���Yof(0=�����K�he��?��=�����Hbo�ݖeA�؈�?r���u5�C>>��A�A��������C@#�����>�>>@�����E�A�i�>ښm���+?n0g�y"ϝ n��P2��žR?�?�����J�=� ߿?T-�^���A����<��G���%@��"�j�+�.���CAҙ�����B�r�4�Z�׋ޞ��*�y»"VBţ��B��%���@a>#������� 7�=;�=���5@,?f�����f;�=f���f>@1��A��t����F=@�
��o�� �ϕ�����5$B�te�����ב��.x�q�¢=B�G��B�����������JOGGGING����7�Z�U�^���8?h���s�<̾��>��s���2n�ecA��&AX����6Z�`0�W���A�)���D�~B�����w�ι�7^�P �Z4�A�	��@�1���+�]���Ϟ�5�kg�9��&{�
s	��o��@|�j/=�ք��$~A��(�>��A/�V!@�ۦ^�����%��3�;��G�$AD?��B�x^���@��?�Y����_�A$F@�x!+�=���U��oJ־�s���)迂������G��נ����@� ����,A�7A���BP����N�Js2��@����l2B��wy��E����ҸN<��������'�7����¤ǌA��Y>:��@��oJB�;ż�V]�/d��@Sp[?���@,������^�w����)A��A�m��Bi�������� �@�����k�����տD���ѩN�� �����~��G�¬�tOA��7#5OB��LO�{�����
G@�w�?p��i?�¾r��17^����"���A���Ae�ӴA��-���T�?@����ԳB�i���Z/�����N&����v�h�O?���ªX�A� �P�	�Yq�U<�XX�=��=���;Y�3<ӕ:+NN�h���3�A���@��T��8߬�WSQg>�B�A��������B�Ę�֌���Ԙ^��� ?����AY�A�D�4��7@@g����5NL��ML�U��4p��tey=L��>6�T�R��>�Ύ>?����j lA�m�@��ɿP�O�j
nB�b����^���n�B����֞`����)7^���!��jA]�3AN�g���/@ s���̚@PAL�/��=!VtzڛU>�.~����������-w?G��?{W�N��`����AΥu�sq@���-#�����qA�L���HƉBO�Al�Cp\�o`F"kAC��ƿ �AG��>����W�ASSEMBLY ER�?�.�tz�6�+����;��Cj�>��^=�%��1�o��'ݰ���Ȁ'��PK_@�X�@�`�?�EA���I�B ���Alc>C���7��B`�T���!�1A-?����)mGOYO~>_ VA`��U�?!;��
���I�>��Z���Wh���$�/�2��[�	�AЃ�?!���@��@8����W�4AV�y��T�N�B�*B�qFJ��,@��,��A5�A7xw�@�<�}�2M�ASTER��j�VAb���:a���>�ڴ@ϖ�� �����L�^��ڼ�A�[�?��Ah�>p?D�v���]`a-A~b�6�Ң�~`�C4y뿢�����q��-O�Z��mA+)@�H��O�DOOR ���6_�g'`�WV�����1���Y��S?��C���&�y�ߞY�N��9<A��}�?`�>AC�T�?�\	�Q��XA�Q}���s�J�BM�l�CY��~�����(IA��f@ԿoA&��w��[�ok�6^���&{;c6��:�W~��=����w-=���v�ۍP���(��@�@�A�=fso]`_���A����  �B�N�UP	�hTAR��?����A��!���bO�=�2Q�����VAs��6�8(�@�>��S�@j��w;w��8��T�W���LA��#?���A3Z@�g%2{����,]A��B��,�`�YB�N��/��e�7��b�UU@�@�!d=�]\�]�d��VBdi��=$��w��;^���nl�W�,@�%�A���������A���h@�G�@s�s���/���>V�8E�A(�U�A���ʿ� ����ۮ����n�e@k�����A=��C�cEOg�4��w����&ڲ�@Ӝ��?J�A5��ʿ��*�cl�������)�jA�u�?�j�a>��h@���
[ΌnZ����
�{VdB�V���Rt�̣��[έE����4Ake�A����r:">�h�c?�=�*�h���%���F��j4��N�S��o߿BJH?<ww-�����A��.@��.����������Y���!�����B�m��ϟs���d���Q��n@�c�@��~���,�%p�\ ����Bd����>�25�?��B���/�vU��	��H �A�g�ῇX��@*��^p��Aλ��p���B����G�������d��8@���@���@�����:���^ ��ϴ�7�����=��?�����>X�ܽġ/��6^*�=T��0�AՑU?VrS��&��@[�I�?�f�Aص����>B����k�W��-E&�A�-s�@�i��:`�O��Ϭ�φ� 6���%���དྷ��=�!���k=����=�tV��<���X4PA��@���x�]M���N�n9A�*�����B�WS����s���ǎ�G������A���@�����$	?����|TTAU�eQ�\��
VBeӟ�;	����w�l:�?������}c���>��$lA���?d�7�?��?�4�K��3<A�q����sB������T�����P��&��A}�A� �h���A���mp�)�D�e�+i��з>�!����>	z>���<��z�Aם����(��)�����3�A�c�U�X%�B����ܳ�����w^�%%��S�iA���@1�yG 6�:�������fN�y<�=H?��g�:���#/Yd0��A���>��A�ߐ@&�w-�	��8�n�@���(��`����B���C��PAt��[A�!�?�V�AP����kb
��a�?�*Bh�&@6�lA���A��@6���{��1�-��������A��%?����AU[@4+��N:-�������7 �Bq�CoϢ��(Ԍ�'�_�A� �A��@�%�?DO������}o� 2�����A�������?�нAt�?�,^�}��A�h!A.��c��(����#>%��BJ������OB�5�}�+@�A��Xg��8��!�A{S�@w�e�� �@Q�pJ��4U�/�,$���+f��?$] @�z������e?���_��h�����A��ӐA??������N"�Q�X?�CB�����(ff?��8�o���@3��A�@���m@�*H@\��[/m/R?� NV��վ����1�#�>�d�1�����;?����w^�bo���@A��A){������_�A�3A�o���V�RB��m��z�Иx�N��P��0�A,EzA%�|����?�A���ASERM�ARK�(GVN�XZ�fVk���li>[��]���@P�A ����*������
A�A
���@w����w^�F�,���@��B����A5�!�A���Q�T�A��]��)��AC��As)����OI�Nd�#�����E:0 ����=��}�������A��a�+a��@����ǎ�����l�@��+��^R=�!UjC�)�^��|������_�@�1���߰���V��Nv��f���^?\��>@�[F��+����G�?���ǎ9�q�#�(���2�=� �ICm�_�~	����]��͖�����CC ى�>�P�5QоC����	r�p95��>Q�S O]��VNz��f�c�A�"A!��>�s?����>
�ǎ?����ĊA���@������<￿���>�f��A:���z�B�W����x��o�����XA�2��AfPj�((\��'��Q�i��N���g���=J���2Y��?K���t@���` �h���A�Q�A/��a@�p��u5�_C)����El���s±���B���B��c�>��@��0�@��Ao���?xa���/?CONVEYORSֿ�L��p�չ���m3Ύ�;��{d;,PAB��>���L��t�A��q{��Ơ@�����Z�r����_�A�����GK��� ��Z_�\�����A}��?�j7�A�eLA�,=L��o�N�j6@�&l�d>��K@͏�٫[��ks���p�T�A�w?�@c�9@�V��@����~$�b��0�?�_3�¡��B�v��B�,����_Z A�ұA�ݠ8,4�V�'��9��U��#�&�k�)X�������g=Zzߙ>��];�5���j-���@������T��~���A�����i9¥�B����B�I�J����B`�k0+@���A�A@R�2s���D���h�O�KY#�ԏ�� ������N������@��;ހA���A�Ň5@3J�Ab|�p�/n�]��@���A1����?�)bίO��A��AV(�?����A-��?�n0�OASSE�MBLYȯ��	V�O���9@��RZ���-?��0@F��?��B�;�<����^��A��@���C�԰W������.�@v��	m;�.�EB�����ՙ�C�*�O���Z4��@nYAh���@~=���� ��>3F2I?p���b��������S��\2?.����v͚?�>(�;�J$l�D5��A��@z{�?���N�B���������S�r5B�f3�߿��C%åO�����0@MOK�Au��0��5!:ZZW�<�D�(��F���>��@q���@-��D��>�tA���_Oq@��A��%�Am������tBX=�.��Zk��Y����B����?�tC)giO�����\x@�@0@�d\�A��#���e�1�� +����[�!t?t�A�}1������>P}ƿ^�n{�q@��sA����A�m���gmBȦ�B��r���%���JGB�c�����p�M��1��P�(��@�J��?��dB?��Ƌ/��������c�s�,.�,?�s?-��%=���?9e��Tn�nZ��J���AdI���1�@j��+@X_�Q���mI�A�����r���±�B��"����:��Y-
A�I����A��_?�����er�����VO���u���?^sY>����>�y>�o��Y�5[^L��f�Ț�A��X#�@��@B�;|/n�ӿ��{��~r�A���zA�L�Bm�z�����wA��
���A���Yyɛ��eq�ET���
�VO��c�>�$�;?��������+��?� �0@���[^E��u��UA�0@�k�)@�1�N��_����Sx�'@��C�t���**�r��9?���b�:�AB���N�q�A|<�@�vy�o�f���c�����_��͹?�
:?wvy>�������������y�LA����;�	�A*�*�Х��/��>+�CUA0�b �CZN[^�S���яA�wQ��p��3+ ����:_x���-O��'< ������>8I�>��O:=��H����������u���A��A3�4�c�@����������E&��CTKM�h��C."�3^�����A�����V��L1����K/��?M"[��_9�&{�;�:����:�=���p�3^TP���xA����F�s��`�A�F>���C���F���CTf�i�V��������=�E�A"���?d �#P��� ^J�/�?G(��c���m32���w�?2��q�ͽ�(`���,A�5��D�v��c�5A)/.o?�{��0��F���0g>�0{B���ӎ<q��BI@�&������T��Fal�?�?�OM!�{c���7u��o��
J���t����B�?i�E��Ϲ��q��x@חSQ>��<�N_����6�����^B�K������ҏ:����;^AU�U@����"&��=����LEAK�TEST ��W�VO�c�o�k����w�l��W�~��A�0���6�Β����A��@�@������ H�X�������->���*B�h�$�̽�D�G�>v����r�A��w@�����?,4@��7�Oer��@�`h*�Pc�;�� �=��W��eˉA*F������Q?�>�'ݰ��NA��@�t�A!��A�C�_��������JE�B:M4�7l[������|������@��R�@�"@�.�� �vg_yV)�����a��<�j�N��=���;ӕ�V�hw{�`�>����C�?D��?%�:��o���,_���+�`]`ߧB�������T�AH��AZ��@. � '�;o�&�do��9<&{��^�>�LJ�F1�`tVN�P���Aǹ��?������h@)���4���+���-��B�|�$���B��������AR�����25?�)m�!ڏEr��Fɏ���W%����@ƽ��~&�����{\	��>��Aم͞c�@�7���������:����Q�B�ܝCrũ�>�d����MA)�RPA.3@�?$�?c�뷏y_쮟�Q�wf����=����\ox�A*����߇��0�W��R�Z���v�A�H}��VrS?�Β�@�5g�"����gi��SB��]���������&����A �AF�����:����߰��������S���:����40>?�G�::І�����}p�Y�A��5�@�?ط�?�� ���� ������$ѵE��B"%Cu1�rk~��>Ş�A��@�@�@߹,q��,J?OGGINGy�/ �z�Y����������m� |���5:mW~9���=��6�>}��}�A�m�C@�&v@������b����m��	P �1B��Cu �s.�
��ah��A��A4@�0��e\�@�!�`�PGH�Y?��Ѕ?�(9񞱯��̡��:A���@��牋mO������)���!�`}^`F���>�-%�cA���@�����6?���E���=��I�(�>����h`�����A6&A��;o վ�����A�b�@����@@y����s.�������J��˧AD3��@��B�i��s.�����W@Ց��%�*A�f�AS�����B��Uo��3V�PK���?�������<�ˉ���
?����@�R�kN�)���p�A�D��@��*@u5���ۦ�n���[^A����@\=:��&@�B���n�▇����,A/8���J��~=@��.eCU�� V�PR��������~�?������M���A�1рo�����A���@���AC�x��p�CN����W���A�*@A��/�����B~��js.1�P���Q����V�AX3�A4� �ڝ��S L��|�
����F;dg�����w�t@^�����/G>`���[��A؈��_<B����{@tT�CNw� � ����Q�"C1�`��ج³H��kN�E���ާ�O��2�ߦ�\͒W�S �PV�PW�F��
���ȿ��@��E��s֋��t�.��X����	�A�&����ݰ�L�f@��U[CN?�|��;u�J��CG�q4�D/k�����>3�����)A3��?�������俛�V��ߥO" @V�P]�V?�q�@���@��@�(�@SQ������J�����eA����|�=?�ք@a��<c���~��z���eHnA��$A��5B�r�2���q�3��A��濯���A����ns0�BLY$��M�P.�$SE�RV_MAIL + _�% ��$�OUTPUD &�3$RV� 2g�  (  (�TJ!�P�Rx(<�$SAVE;,))�TOP10 2�[) d �� �R��2�Ps��s*�PO��r�Pc��/ ??1?C?U?g?y?�? �?�?�?�?�?�?	OO -O?OQOcOuO�O�O�O �O�O�O�O__)_;_ M___q_�_�_�_�_�_��_�%YP�/+#FZN_CFG �(#�J!�%a�GRP 2����! ,B   �A_`�D;� B}``�  B4]ÿRB21�&H7ELLbcŪ&�z �. 6g�o�k%RS���o�o" F1jU�y�� �����0�B�T���  �c!%@U�����c�����K 1������ޚ�k���!d�����fHK ;1�k ŏI� D�V�h���������ٟ ԟ���!��.�@�i��d�v����lOMM ��oد�bFTOV_ENB$c!�)�HOW_REG_�UI��,"IMIO/FWDLàǮbe^-�WAIT�����7bU�5 �b$R�T�I
 �����V�A c�-�_UNI�T��ö�)LC�T�R���% M�B_HDDN 2[+ 6���>� 4�`�U�h�P�bϏφπ���ϼ�������O�N_ALIAS y?��F#( heb! 7�I�[�m�߉�3߬� �����ߍ���*�<� N���r�����e� ������&���J�\� n���+����������� ��"4FX| ����o�� 0�Tfx�5 ������/,/ >/P/b//�/�/�/�/ �/y/�/??(?�/9? ^?p?�?�???�?�?�? �? O�?$O6OHOZOlO O�O�O�O�O�O�O�O _ _2_�OV_h_z_�_ �_I_�_�_�_�_
o�_ .o@oRodovo!o�o�o �o�o{o�o*< �o`r���S� �����8�J�\� n���+�����ȏڏ�� ���"�4�F��j�|� ������]�֟���� �ɟB�T�f�x�#��� ����ү䯏���,� >�P���t��������� g�����(�ӿL� ^�pς�-Ϧϸ����� �ϙ��$�6�H�Z����$SMON_D�EFPROG �&������ &*SY�STEM*aߥ��@�s�RECA�LL ?}�� ( �}�����&�8�J� ��o��� �����\������#� 5�G���k�}������� ��X�����1C ��gy����T ��	-?�c u����P�� //)/;/�L/q/�/ �/�/�/�/^/�/?? %?7?I?�/m??�?�? �?�?Z?�?�?O!O3O EO�?iO{O�O�O�O�O VO�O�O__/_A_�O e_w_�_�_�_�_R_�_ �_oo+o=o�_aoso �o�o�o�oNo�o�o '9K�oo�� ���\���#� 5�G��k�}������� ŏX������1�C� ֏g�y���������T� ���	��-�?�ҟc� u���������P��� ��)�;�ίL�q��� ������˿^���� %�7�I�ܿm�ϑϣ� ����Z������!�3� E���i�{ߍߟ߱��� V�������/�A��� e�w�����R��� ����+�=���a�s� ��������N����� '9K��o�� ���\��# 5G�k}�����X�$SNPX�_ASG 2������� P 0 '�%R[1]@g1.1�)?�X9%/B/ �(/i/�t''/�/�'��@�/�/|/�/�/Z��/'?38�?Y?c6G��H?�?�6�?�?J*ܨ?�?�/�?OZrVOIO�?>OObO�OF.j�O�OL(���O	_�O�O?_Z��(_i__^_�_�_ �_�_�_�_f�_'o�_o]oYoFo�o:o |o�o�o�o�o�o�o�M0q�~�� h�\�������9��.�o�"�����MN��ɏ�? ����R�#���Y�d��+H�����BC8x���Ö�G��� ̟ޟ�B�C���8�y������h�����I ��ׯ*�̯��1�C� �(�i�/^���R�ÿ տ�������/��S�0�Hωϔ�
�xϹ� <Ϯ������%��I�p,�>��ZP 1h� ��\ߞ��������� 9��.�o�R���� ���������)���`�_�B���w� x�������������B����l�OZ2 ��w��h�,�����PARAM ��� ��	_P��S!��=�t��OFT_KB_CFG$��p���OPIN_�SIM  ��2���T � RV�NORDY_DO�  <h�QSTP_DSB|�2/�SSR � � &� PNS001�0 MBLY D� /�n�OTOP_?ON_ERR��~�!PTN �� �C�"RING_PRM�/��VCNT_GP� 2 @Bx 	/?1@�/6?!?�Z?+'VD� R��!AK17E7�?�? �?�?�?OOO%O7O IO[OmOO�O�O�O�O �O�O�O_!_3_E_W_ i_�_�_�_�_�_�_�_ �_oo/oVoSoeowo �o�o�o�o�o�o�o +=Oas�� �������'� 9�K�]�o��������� ɏۏ����#�5�G� n�k�}�������şן ����4�1�C�U�g� y���������ӯ���� 	��-�?�Q�c�u��� ������Ͽ���� )�;�M�_φσϕϧ� ����������%�L� I�[�m�ߑߣߵ��� ������!�3�E�W��i�s2PRG_CO7UNT]�"��'ENB�/��M��_���_UPD 1">:+T  
~�& �#�5�^�Y�k�}��� ������������6 1CU~y��� ���	-V Qcu����� ��/./)/;/M/v/ q/�/�/�/�/�/�/? ??%?N?I?[?m?�? �?�?�?�?�?�?�?&O !O3OEOnOiO{O�O�O �O�O�O�O�O__F_ A_S_e_�_�_�_�_�_ �_�_�_oo+o=ofo�aoso�o�o�o�o��_INFO 1#�����p	 ��o"F1y<���<3���ft�;fpQ}B�����`d�A�BN;�:�����wB����Q}?�@ �D��C�9���aACPL ��7 D���D���B���8�|y�  ���w��YSDEBSUG�� ���`d����SP_PASS��B?"�LOG� $�f	�  ��`h�?�ה��`�o  ����a?UD1:\N��n�O�_MPCT� P����ۏ����2��~��SAV %W����8qw�׊��S�V�TEM_TI_ME 1&W�
� 0 )��ck|��� ^�c��`�MEMBK'  ����w�w������X��'� @����(�M��]�!�������� 8{@��į֯��� 4��%�7�I�[�m�� �������ɿۿ� ���#�5�o�eD�i� {ύϟϱ��������� ��/�A�S�e�w߉�0�߭߿�b�SK����@��ϟ���#���P�p%�	�:�j��` �dáo����N 8���������8}� �0�  �W��i�{�����������������
.�`A$2VJ�z�d{� ����� $ 6HZl~�������gT1SVG�UNSPD8� '�"���2MOD�E_LIM '�t�&��2�!(�W��ASK_OP�TION�Ù&��Y!_DI1�ENB�  ��"�y!BC�2_GRP 2)���"����/j���C���#�BCCFG +�+Ս.�׏:`$?S\?G?l?�? }?�?�?�?�?�?�?"O OOXOCO|OgO�O�O �O�O�O�O�O_	_B_@-_f_Q_�_�_�d�\ �_�_�_�_v_�_1oo Uo@oyo�j�՝oɐn` �o�o�o�o�o�o3 !CEW�{�� ����	�/��S� A�w�e����������� ��ۈ�P	��9�K�]� ۏ��o�������۟� ��͟#��G�5�k�Y� {�}���ů���ׯ� ��1��A�g�U���y� ����ӿ������-� �Q��i�{ϙϫϽ� ;���������;�M� _�-߃�qߧߕ��߹� ������%��I�7�m� [����������� ���3�!�C�E�W��� {���g������� ��A/Qwe�� �����+ ;=O�s��� ���/'//K/9/ o/]/�/�/�/�/�/�/ �/?��)?;?Y?k?}? �/�?�?�?�?�?�?O O�?CO1OgOUO�OyO �O�O�O�O�O	_�O-_ _Q_?_a_�_u_�_�_ �_�_�_�_oooMo ;oqo'?�o�o�o�o�o [o�o7%[m M������ ���E�3�i�W��� {��������Տ��� /��S�A�c�e�w��� ��џ�o����+�=� ��a�O�q�������ͯ ߯����'��K�9� [�]�o�����ɿ��� ۿ���!�G�5�k�Y� ��}ϳϡ�������� ��1��I�[�yߋߝ� ��߯����������9��$TBCSG_GRP 2,���  ��9� 
 ?�  d�v�`����������������(�=�D�.K�d���Y�?9�	 �HC� (�&fafu�9�(�i�A�9ἒ���D)�(�c�ͽ�)���B4�������L��~�����/Cj����3�33(�B�C/1C(�a��f)�>����Bܿ@~��~�-@ k�Se�������	V3.�00�	rc2l�	* $8��*/�G�?�3e39�XM!� a 3-b/  ���/��%=�J2D�/K���/�(CFG 1��U�]��*��\�w"�/68�6?\?j:�j?�?{? �?�?�?�?�?�? OO OVOAOzOeO�O�O�O �O�O�O�O__@_+_ d_O_�_s_�_�_�_�_ �_oobv�#o5oGo �_zoeo�o�o�o�o�o �o�o.@Rv a����9�%�� ����O�=�s�a� ��������ˏ�ߏ� �9�'�]�K�m�o��� ����۟ɟ���#�� 3�Y�G�}�k�����s� ˯ݯ������C�1� g�U���y�����ӿ� ������	�?�-�c�u� �ϙ�SϽϫ������� ���;�)�_�M߃�q� �ߕ߷��������%� �I�7�Y�[�m��� �����������E� �]�o���+������� ������/Se w�G����� +�;aO� s������� '//K/9/o/]/�/�/ �/�/�/�/�/?�/5? #?E?G?Y?�?}?�?�? �?�?��OO�?�?UO COyOgO�O�O�O�O�O �O	__�O+_Q_?_u_ c_�_�_�_�_�_�_�_ oo'oMo;oqo_o�o �o�o�o�o�o�o 7%[Im�� �����!��1� 3�E�{��?������a� �Տ����A�/�e� S���������}��џ ����=�O�a��-� ��������߯ͯ�� �9�'�]�K���o��� ������ɿ���#�� G�5�k�Y�{ϡϏ��� ��������ɏ7�I� Ϗߋ�y߯ߝ����� ��	���-�?�Q��!� ��u���������� ��)��9�;�M���q� ��������������% I7m[�� �����3! WEg�{�+�]� ����//S/A/ w/e/�/�/�/�/�/�/ �/??)?+?=?s?�? �?�?c?�?�?�?�?O O%O'O9OoO]O�O�O �O�O�O�O�O_�O5_ #_Y_G_}_k_�_�_�_ �_�_�_�_ooCoUo �moo�o;o�o�o�o �o�o�o	?-cu ��W�������~  +�/� �/�C�/��$TB�JOP_GRP �22�u��  ?�/�	�[�b�4i���p� �� ��,^~� ��� � s �� �/� @�+�z�	 �C�� ߆Qp�D�q�/�z���&ff�x����<9]߁�?��?L��~7�BH  A���<R�]�D)�o���S�Y9����� ;�<�>����<��o�?33�3?f�ȐB� � B I��m�D5m󎴔�$�8�8��,�Af�ÒD�{�C�ؐӑ۟|�Cj�����|�.�ȑ��ª;�?��B�ǖ���a�}�
�����1��<�N�<��㪌��󯔿�)��������ϿՀ̑̐��z��J�|�>���C4Ր���*�ɿo�C� ]�G�yσϴϏϡ��� ����	��D��1�c�@}�gߙߣ��ߧ��/�������	V3.�00��rc2l�*!��*�/�:�� F�  F��  GX G�7� GR� G�r0 G�� G��@ G�� G��\ G�� G��` G�� H�
� Hd H�" H.� H�;� HH2 H�U�J�E�� E|T��F@ F���Fj` F�� �F� O�|��� G$ G��G�V�b㈸ G��L G�� G��h G�� =u�=+��X��k�9��1�5�?�  Ӆ��M��ESTPAR°�#�t�X�HR��AB�LE 15i� IS�/�:船)�
:�:�:�.�6�:�	:�
:�:���/�U:�:�:���'RDI��s����� �����O��@�������S�q� O
����� //0/B/T/f/x/�/ �/�/�/�/�/�/?N� ��r���I92DV h&8J\n��~/2NUM  �u�s�π7� ���� ��_CFG �6K�3Ӂ@[�IMEBF_TT��p�5q���ZFVER~�[1pFZCR 17��� 8,�/�d*��A �pT?  �O �O�O�O�O_!_3_E_ W_i_{_�_�_�_�_�_ �_�_Boo/oxoSoeop{o�o�o�nDAC�o�o�n	$B�o�n�_TM1C�nT3�oz� ؒ����jILL���~Pc_A�#��~$M�oZ�l�ER�@����L=# ��ˏ�D_A�F�@�E��MI_CWHANfG �E 4��DBGLV�hE��E��7�ETHER_AD ?����m�5�0��:e���4:79:ee:�f5 ��6��f7���f8q�ROUT6�@!!���~�7�SNMASK���C��255.E��C�U�g����OOLOFS_D�I°�i�ORQCTRL 8�K�6��Tԯ	��-� ?�Q�c�u��������� Ͽ����)�9�ӯ�\�Kπτ�PE_D�ETAI]���PG�L_CONFIG� >I(A���/cell/$C�ID$/grp1�������0�B��� �om�ߑߣߵ���V� �����!�3�E���i� {������R�d��� ��/�A�S���w��� ��������`��� +=O����������S>}t' 9K]o�1qϗv�s���//&/ mJ/\/n/�/�/�/3/ �/�/�/�/?"?4?�/ X?j?|?�?�?�?A?�? �?�?OO0O�?TOfO xO�O�O�O�OOO�O�O __,_>_�Ob_t_�_ �_�_�_K_�_�_oo (o:oLo�_po�o�o�o �o�oYo�o $6 H�ol~���������User View ���}}1234567890	��-�?��Q�c�k���Ë����y2�yh͏ߏ�� �'������r3��u� ��������ϟ.�🞎4d�)�;�M�_�q���⟤���5�ݯ��@�%�7���X���6̯ ������ǿٿ�J����7��E�W�i�{ύ������Ϟ�84���߀�/�A�S߲�t�z� �lCamera�z�Ϲ����������E��=�O� a��{��������˩  �֯���%�7� I�[�m��&������ �����!3El����c������� ����!3~W i{���Xj� H�/!/3/E/W/� {/�/�/��/�/�/�/ ??�j��/k?}? �?�?�?�?l/�?�?O X?1OCOUOgOyO�O2? ��� O�O�O�O__ /_�?S_e_w_�O�_�_ �_�_�_�_�Oj3Ɍ_ AoSoeowo�o�oB_�o �o�o.o+=O aoj���o��� ����o+�=�O�� s���������͏t�w9Y�� �2�D�V�h� �y�����W�������
��.�@���	��0 Ɵ{�������ïկ|� ����ğA�S�e�w� ����B�T��М�?��� ��*�<�N���rτ� ��Ὼ��������� �������`�r߄ߖ� �ߺ�a������M�&� 8�J�\�n��'�a�t ���������&��� J�\�n���������� ����������8J \n��9���� %�"4FX�� ��L;������ ��"/4/F/�j/|/ �/�/�/�/k��K[/ ?"?4?F?X?j?/�? �?�?�/�?�?�?OO<0O�-  �)_O qO�O�O�O�O�O�O�Ox__%[   5O =O[_m__�_�_�_�_ �_�_�_o!o3oEoWo io{o�o�o�o�o�o�o �o/ASew �������� �+�=�O�a�s������)\  
� (  ��S@( 	  ��ݏˏ��%��I� 7�Y�[�m�����ǟ��t럱�EZ �? 0�B�T��?x������� ��ү�#���� �g� D�V�h�z������¿ Կ�-�
��.�@�R� dϫ��ϚϬ������ ����*�qσ�`�r� ���Ϩߺ�������� I�&�8�J��n��� �����������W� 4�F�X�j�|������� ������/�0B Tf�������� ��,sPb t������� 9K(/:/L/�p/�/ �/�/�/�//�/ ?? Y/6?H?Z?l?~?�?�/ �?�?�??�?O O2O DOVO�?�?�O�O�O�? �O�O�O
__._uOR_ d_v_�O�_�_�_�_�_ �_;_o*o<o�_`oro��o�o�o�oo�@ A�b�o�o�c�g�ǀ��)frh:�\tpgl\ro�bots\r20�00icGu_12?5l.xml�oq �������������D�V�h� z�������ԏ��� 
�!��@�R�d�v��� ������П����� �<�N�`�r������� ��̯ޯ����8� J�\�n���������ȿ ڿ�����4�F�X� j�|ώϠϲ������� ����0�B�T�f�x� �ߜ߮���������� �,�>�P�b�t�����������&x�\a �o1p<<w /p ?�� G��?�a���u����� ����������C) Ky_�������f`(�$T�PGL_OUTP�UT Aaa;" 7L ^p������ � //$/6/H/Z/l/ ~/�/�/�/�/�/�/7�'��� 2345678901?!?3? E?W?i?q3b?�?�? �?�?�?�?�?�?(O:O LO^OpOO~O�O�O�O�O�O�O�}�O&_8_ J_\_n___�_�_�_ �_�_�_�_o4oFoXo jo|oo�o�o�o�o�o �o�o�o0BTfx �"������ ��>�P�b�t���� 0���Ώ������� $�L�^�p�����,��� ʟܟ� ������H� Z�l�~�����:���د����� ��M'�$$��/b�P���t� ����ʿ������ 6�(�Z�L�~�pϢϔ� �ϸ������ �2�$�V�H�z�}"�ߦ߸���������@)�#�5��/� ( 	  |�j�X��|����� ��������0��T�B� x�f������������� ��>,NPb���6�  <<o��< �*<`r�*� ��O����!/ 3/�7/i//U/�/�/ �/�/�/E/�/?�/	? S?e???�?�?�/�?�? �?}?OO�?%OOO�? �?�O�O1O�O�O�O�O __sO9_K_�O7_�_ [_m_�_�_'_�_�_�_ �_5oGo!oko}o�_eo �o�o_o�o�o�o1 �ogy��� ��CU�-��9� c�=�O�����	���� {�͏�)��M�_��� G���/���˟ݟ��� �q���I�[������ k���ǯ%�7������ �E��1�{���믱� ÿ]�����ӿ�/�A���)WGL1.�XML��v��$T�POFF_LIM� � ������N_SV�� � ���P_M�ON B�Ԡ���2��ST�RTCHK C�����߇�VTCOMPAT��=Ѣ��VWVAR Dr��`ط� ߩ x������_�DEFPROG �%�%PN�S0010��{�_DISPLAY���ި�INST_M�SK  �� ~��INUSER3����LCK<��QU?ICKMEN`���oSCRE��~>�tpsc�Ԡ<����°�_��S�T1ڞ�RACE_�CFG E���`���	��
?�~��HNL 2F��� �g� ��S�e�w����������������I�TEM 2G?�� �%$1234?567890&8  =<0Vhp�  !v~�� :���$�H ~0��}��� ��TDVh�� /�\/�/�/��// ./@/�/d/?6?H?�/ T?�/�/�/x?�?*?�? �?`?O�?�?_O�?zO �?�O�OO�O8O�O_ nO._�O>_d_v_�O�_ �O_"_�_F_�_o*o �_No�_�_�_Zoroo �o�oBo�ofoxoA�o \�o���o�, �P�t �F��� ����~�(�ԏ�� �p�0�������2�܏ ������$�̟H�Z�l� �>���b�t�؟���� �ׯ2��V��(��� >������毦�
��� ܿ�R���v������ ��jϐϢ����*�<� N����τ�D�Vߺ�b� ���Ϲ����8���
�@n� �ߤ�m���S��H�r��  ���r� �����
� ������ ����UD1:\-������R_GRP 1�I� 	 @��x���t�������������� '
���-�Q<u`?�  ������ �
�.dR �v�����/�	@�/,/��SC�B 2J��  {x/�/�/�/�/�/�/��/?x�UTORIAL K���S?�}�V_CONFIG L���o�����?c<OUTPU�T M��0���?OO&O8OJO \OnO�O�O�O�O�O�O �1�?__&_8_J_\_ n_�_�_�_�_�_�_�O �_o"o4oFoXojo|o �o�o�o�o�o�_�o 0BTfx�� �����o��,� >�P�b�t��������� Ώ�����(�:�L� ^�p���������ʟܟ � ��$�6�H�Z�l� ~�������Ưد��� � �2�D�V�h�z��� ����¿Կ���
�� .�@�R�d�vψϚϬ� ���������*�<� N�`�r߄ߖߨߺ��� ���ߌ2��?+�=�O� a�s��������� �����'�9�K�]�o� ���������������� �"�5GYk}� ������ 1CUgy��� ����	/-/?/ Q/c/u/�/�/�/�/�/ �/�/?/(/;?M?_? q?�?�?�?�?�?�?�? OO$?7OIO[OmOO �O�O�O�O�O�O�O_  O3_E_W_i_{_�_�_ �_�_�_�_�_o_._ AoSoeowo�o�o�o�o �o�o�o*o=O as���������������7�I�3�"�t� ����Ώ�����(� :�L�^�p�#������ ʟܟ� ��$�6�H� Z�l�~�������Ưد ���� �2�D�V�h� z�������¿Կ��� 
��.�@�R�d�vχ� �ϬϾ��������� *�<�N�`�r߄ߕϨ� ����������&�8� J�\�n��ߤ���� �������"�4�F�X� j�|������������ ��0BTfx �������� ,>Pbt�� �����//(/�:/L/^/p/�/�+�$�TX_SCREE�N 1NK��3��}ip�nl/� gen.htm�/�/�/??�,?��Panel setup0<}�0?q?�?�?�?�?�?_?U?OO&O8O JO\O�?�O�?�O�O�O �O�O�OuO�O4_F_X_ j_|_�__3_)_�_�_ �_oo0o�_To�_xo �o�o�o�o�oIo[o ,>Pb�o�o ������{(� �L�^�p����������.UALRM_M_SG ?�)��  ������<�/� `�S���w�������ޟ�џ���&�څSEV7  �X�؂ECFG P�%��!  �@�  A��   �Bț� |���{�{�A�;T�̭ϟ�{�@�?v�T�ID��֢@���Uuwz��ѯ���z�A^�Uvc ��a�����iUw����%K�]�o�}�d�GR�P 2Qn� 0����	 @
���z5�>������?���-�I_BBL_N�OTE Rn�T��l�� �z�ڲDEF�PRO�%� �(%PNS00�5��:ϔ%FL?AGSSETE�K� ���|ϵϠ����������!�3��W�շFK�EYDATA 1yS�)��p }�����߼��ߥ��ߌ���,(�2�(�POINT  �]:�<�  OOK� T����i�NDI�REC`ϓ�  C�HOICEU��TOUCHUP�����y�RE INFO��V�h�O���s� ����������
�@'dv ���/frh/gu�i/whitehome.pngw`�������point�1C�Ugy  �look ���������indirec;/M/_/q/|�/�choic��./�/�/�/�/?��touchup�+/C?U?g?y?�?
>�arwrg*/�? �?�?�?O�(*O<ONO `OrO�O�O%O�O�O�O �O__�O8_J_\_n_ �_�_!_�_�_�_�_�_ o"o�_FoXojo|o�o �o/o�o�o�o�o �oBTfx��� ������"�4� ;X�j�|�������A� ֏�����0���B� f�x���������O�� ����,�>�͟b�t� ��������K�ί�� �(�:�L�ۯp����� ����ʿY�� ��$� 6�H�׿Z�~ϐϢϴ� ����g���� �2�D� V���zߌߞ߰����� c���
��.�@�R�d� �߈��������}-���� ��)�@;���d�v��,\���TPOINT� 31��L 1842�� [$H�/TOUCHUPZ[����� ��(L^E��i�����{�"6whitehom�#/&/8/J/\/k�="6poin�?�/��/�/�/�/s�5look�/$?6?H?Z?l? s�?�?�?�?�?�?y? O O2ODOVOhOzO}!��&touchup?�O�O�O�O�Oz$}�&arwrg�/ 5_G_Y_k_}_O�_�_ �_�_�_�_�_o1oCo Uogoyo�oo�o�o�o �o�o	�o-?Qc u������ ���;�M�_�q��� ��$���ˏݏ��� ���I�[�m������ ��ǟٟ����!��� E�W�i�{�������@� կ�����/���S� e�w�������<�ѿ� ����+�=�̿a�s� �ϗϩϻ�J������ �'�9���]�o߁ߓ� �߷���X������#� 5�G���k�}���� ��T�������1�C� U���y����������� b���	-?Q�-_��_�@������,�<�OINTD��hO�s[C?HOICE]�t OUCHUP� ��//>/%/b/t/ [/�//�/�/�/�/�/�?(??L?+�Vw�hitehome %_�?�?�?�?�?��Upoin$_O"O4O FOXO��|O�O�O�O�O �OeO�O__0_B_T_�f_�An6choic?�_�_�_�_�_�?�/touchup��_#o5oGoYoko�>arwrg�?�o�o�o �o�o�O#5GY k�o������ ���1�C�U�g�y� �������ӏ����� �-�?�Q�c�u���� ����ϟ�����)� ;�M�_�q���Z? ��� ˯ݯ����7�I� [�m���� ���ǿٿ ����!ϰ�E�W�i� {ύϟ�.��������� �߬�A�S�e�w߉� �߭�<��������� +��O�a�s���� 8���������'�9� ��]�o���������F� ������#5��Y k}����T� �1C�gy�����\<�}�h0����@
/-�>/P/*&,<? �/4?�/�/�/�/�/�/ �/#?5??Y?@?}?�? v?�?�?�?�?�?O�? 1OOUOgONO�OrO�O �O���O�O	__-_?_ Nc_u_�_�_�_�_�_ ^_�_oo)o;oMo�_ qo�o�o�o�o�oZo�o %7I[�o �����h�� !�3�E�W��{����� ��ÏՏ�v���/� A�S�e�􏉟������ џ�r���+�=�O� a�s��������ͯ߯ 񯀯�'�9�K�]�o� ��������ɿۿ��� �O#�5�G�Y�k�}τ� �ϳ���������ߜ� 1�C�U�g�yߋ�߯� ��������	��-�?� Q�c�u���(���� ��������;�M�_� q�����$��������� %��I[m ��2���� !�EWi{�� �@���//// �S/e/w/�/�/�/</ �/�/�/??+?=?��?;�����h?z?�=d?�?�?�6,�O�?�OO�?9O KO2OoOVO�O�O�O�O �O�O�O�O#_
_G_Y_ @_}_d_�_�_�_�_�_ �_�_o1o�Uogoyo �o�o�o�/�o�o�o	 -?�ocu�� ��L����)� ;��_�q��������� ˏZ����%�7�I� ؏m��������ǟV� ����!�3�E�W�� {�������ïկd��� ��/�A�S��w��� ������ѿ�r��� +�=�O�a��ϗϩ� ������n���'�9� K�]�o�Fo�ߥ߷��� �������#�5�G�Y� k�}���������� ����1�C�U�g�y� �������������	 ��-?Qcu� ������) ;M_q��$� ���//�7/I/ [/m//�/ /�/�/�/ �/�/?!?�/E?W?i? {?�?�?.?�?�?�?�? OO�?AOSOeOwO�Oh�O�O���K�������O�O�M�O_0_
V,oa_o �_l_�_�_�_�_�_o o�_9o o]oooVo�o zo�o�o�o�o�o�o 5G.kR���� ������.OC� U�g�y�������>�ӏ ���	��-���Q�c� u�������:�ϟ�� ��)�;�ʟ_�q��� ������H�ݯ��� %�7�Ư[�m������ ��ǿV�����!�3� E�Կi�{ύϟϱ��� R�������/�A�S� ��w߉ߛ߭߿���`� ����+�=�O���s� ���������� �'�9�K�]�d���� ����������|�# 5GYk����� ���x1C Ugy���� ���/-/?/Q/c/ u//�/�/�/�/�/�/ ?�/)?;?M?_?q?�? ?�?�?�?�?�?O�? %O7OIO[OmOO�O O �O�O�O�O�O_�O3_ E_W_i_{_�__�_�_@�_�_�_oo��k��������HoZolmDo�o�ozf, ��o��o�o+ O6s�l��� ����'�9� �]� D���h�������ۏ �����5�G�Y�k�}� ���_��şן���� ���C�U�g�y����� ,���ӯ���	���� ?�Q�c�u�������:� Ͽ����)ϸ�M� _�qσϕϧ�6����� ����%�7���[�m� ߑߣߵ�D������� �!�3���W�i�{�� �����R������� /�A���e�w������� ��N�����+= O&�s����� ���'9K] �������j �/#/5/G/Y/�}/ �/�/�/�/�/�/x/? ?1?C?U?g?�/�?�? �?�?�?�?t?	OO-O ?OQOcOuOO�O�O�O �O�O�O�O_)_;_M_ __q_ _�_�_�_�_�_ �_o�_%o7oIo[omo oo�o�o�o�o�o�o �o!3EWi{��d �{�d ������}����v,��A��e�L� �������������܏ � �=�O�6�s�Z��� ����͟���؟�'� �K�2�o���`���� ɯۯ���#�5�G� Y�k�}������ſ׿ ���Ϝ�1�C�U�g� yϋ�ϯ��������� 	�ߪ�?�Q�c�u߇� ��(߽��������� ��;�M�_�q���� 6���������%��� I�[�m������2��� ������!3��W i{���@�� �/�Sew ��������/ /+/=/Da/s/�/�/ �/�/�/\/�/??'? 9?K?�/o?�?�?�?�? �?X?�?�?O#O5OGO YO�?}O�O�O�O�O�O fO�O__1_C_U_�O y_�_�_�_�_�_�_t_ 	oo-o?oQoco�_�o �o�o�o�o�opo );M_q �� ����~�%�7� I�[�m��������Ǐ�ُ�������>����(�:� L�$�n���Z�,l��� d�՟������/�� S�e�L���p������� �ʯ�� �=�$�a� H�����~�����߿� ��'�9�K�]�o�~� �ϥϷ��������ώ� #�5�G�Y�k�}�ߡ� ���������ߊ��1� C�U�g�y������ ������	���-�?�Q� c�u������������ ����;M_q ��$���� �7I[m� �2����/!/ �E/W/i/{/�/�/./ �/�/�/�/??/?� S?e?w?�?�?�?�/�? �?�?OO+O=O�?aO sO�O�O�O�OJO�O�O __'_9_�O]_o_�_ �_�_�_�_X_�_�_o #o5oGo�_ko}o�o�o �o�oTo�o�o1 CU�oy���� �b�	��-�?�Q� �u���������Ϗ� p���)�;�M�_�� ��������˟ݟl����%�7�I�[�m��$�UI_INUSE�R  ������� � n�r�_MENHIST 1T���  �( ����0/�SOFTPART�/GENLINK�?current�=editpag�e,APP_MA�STERS,1 � ��-�?�Q���+����CUBEIO����������ҿ��'�k���menu�158�3�ST����2�D�V����|�
�P?ALLOAD����������,sυ�PNS0010�2�D�dV��(���07�5,9 �)߽���0��係��74�#� ���@�R�d�����1���0���������������#�5�G�Y�k�}� ����� ���������� 2D Vhz	���� ��
�.@Rd v������ /�*/</N/`/r/�/ �/%/�/�/�/�/?? ��8?J?\?n?�?�?�? �/�?�?�?�?O"O�? FOXOjO|O�O�O/O�O �O�O�O__0_�OT_ f_x_�_�_�_=_�_�_ �_oo,o�_Poboto �o�o�o�oKo�o�o (:%?Cp�� ����o� ��$� 6�H��l�~������� ƏU�׏��� �2�D� V��z�������ԟ c���
��.�@�R�� c���������Я�q� ��*�<�N�`�K�� ������̿޿��� &�8�J�\�n����Ϥ� ���������ύ�"�4� F�X�j�|�ߠ߲��� �����߉��0�B�T� f�x���������� �����,�>�P�b�t����q��$UI_P�ANEDATA �1V������  	��}`/frh/c�gtp/flex�dev.stm?�_width=0�&_height�=10����ice�=TP&_lin�es=3��col�umns=4��f�on��4&_pa�ge=t��1 e�v��o�)pri9m6_  }b�`����� )� �*N`G� k�����//��8/o��� �   h���pa������!2��	2B/=
dual�/�/r#? 5?G?Y?k?}?$/�?�? �?�?�?�?�?O1OO UO<OyO`O�O�O�O�O�F/X" hӲa��h/z/�/P3�/�/#3�O=	thirdv_�_?�_�_ �_�_oo�OBo)ofo xo_o�o�o�o�o�o�o �o>P7t�O�Y! C�a� R������� g8��_\�n������� ���ڏ�ӏ���4� �F�j�Q���u���ğ@���ϟ��Q" �� 8���T�Y�k�}����� ���ׯJ�����1� C�U���y���r����� ӿ�̿	��-��Q� c�Jχ�nϫϽ�0�B� ����)�;�Mߠ�q� 䯕ߧ߹�������� h�%��I�0�m��f� �������������!� 3��W����ύ����� ������:���A Sew���� ��� =O6 sZ������ d�v�49/K/]/o/�/ �/��/*�/�/�/? #?5?�/Y?k?R?�?v? �?�?�?�?�?O�?1O CO*OgONO�O�O/"$��O�O�O�O_#_5_)�OZ_�%I_�_�_�_ �_�_�_G_o�_(oo !o^oEo�oio�o�o�o �o�o �o6�( #�+�$UI_PO�STYPE  � %� 	�p��~hrQUICKMEN  w{���jpREST�ORE 1W %�  ��*defau�lt�+  RIwPLE�}T(��� meditp�age,PNS0072,1�z��������S�menu>[�148,2���p��
����200g� T�f�x����)���� $�֟���#�5�G�� k�}�������V�ׯ� ����ʟ,�>�P�¯ ��������ӿv���	� �-�?�Q���uχϙ� �Ͻ�h�������`�)� ;�M�_�q�ߕߧ߹� ���߀���%�7�I� ����h�z��ߞ����� �������3�E�W�i� {�������������}oSCRE�p?�}u1sc�Wu2(3(4(U5(6(7(8(�TATs}� x�s %`zUSER
 L!ks*�3�U4�5�6�7��8�hpNDO_CFG Xw{�@�A�hpPDk�	�?None�r� �_INFO 2Yj %O�p0%�� j�(X�|��� �/�)//M/_/B/��/�/x/�/�|<OFFSET \wyS�/�����
?? .?@?m?d?v?�?�?�? �/�?�?�?O3O*O<O iO`OrO�O�;��M�O��O
�O_��<W�ORK ]G��O_T_f_�/� UFRAM,�-U9�RTOL_ABRqT�_7�RENB�_~�XGRP 1^�y��qCz  A� .c,a��,o>oPobotoB�f�o�o�Z�pU�X��[MSK  h-UO�[N�Q%G��%�O<�U_EV�N�P�dQv�2�_�+
 h�UEV�P!td�:\event_�user\@�pC�7��O��F%]�pS�P�q�wspot�weld�}!CA6���* +t!+ �m���M��a[���� Տ
���Ǐ@��d�� !�3���W�П{���ß ��<����/���s� ��S�e�ޯ�������ѯJ���n��+�pvWf>P2`�	Q8i�ҿ� ��	����?� Q�,�uχ�bϫϽϘ� �������)��M�_߀:߃ߕ�pߦ�������$VARS_CO�NFI a�+ F�P�����CMRvb2g�+�i��	SR%1:� SC130EFG2 *i�m�����8Y�,��`�5���?�~`@~`p�`�N�� �_���� ������+�P�&�S���-�eA��?�����b B��� ��a��7�������� <'`K]� ��w�����&,8��IA;ThC]/�,		�Au��G�P Ǣ*XN�SIONTMOU�[ ��xri��ᦌ�#a FR:\��\DATA<� � �� MC��LOG/   oUD1�EX'/��a' B@ ��j";!�߈/;!��/�/2� � n6  ���Z��g"�f�'��  =����1a�� < >(TRAINQ/�"42N�dF3p58Da#.T�p�,�j{ (�R9�=�	�? �?�?�?�?OO<O*O�DONO`OrO�O�OIS�_GE�k{�`�`�
(`�R�JN �RE�liSV��L�EX�Dm �H�1-�e?VMPHASOE  uG������RTD_FIL�TER 2n{ Ԋ�ȸ�_�_�_ �_oo)o;oMo_oZ� �_�o�o�o�o�o�o�o�/FSHIF�TMENU 1o}<w,%w/����k���� � ��6���E�~�U��g����������	�LIVE/SNA��%vsfli�vP^���� �SETU��menu5�:�ԏ����|�Ku�pZy�EwMO��q<^�z��ZD�ʔr_<D0�@��$WAITDIN�END�G�ޒ3�OK  C�N��i��S}�P�TIM�����G:�ʭ\���|�ͪ��ͪ��N�RELEgQ��ږ3���{�3�_ACT����dN�_� s�\�%  RIPPERCH����C���RDIS�~���$XVR6Qt~<^�$ZABC+�;1u� ,D0��2�A���VSP�T v<]J�7$
������x���|�ϙ�DCSCH8P�w\��Q�IP�x���ߨߺߓ��MPCF_G 1yr��I�0G�r����MPY�zr�o1��Ƽ���Z�(����  �]���������8BHt���}�?z�dV��7 D��Dׯ��0�A@�
s�z4 >���Q6tT��?�t?��e�w� ���������0)A��_�I����B��8�|y�� ���������������;�������: �#�O���8P{r߮_CYLIND�Q�|�� �0& ,(  * 7#`�:!^E w� �����J�� �5/xY/k/}/��/ </"/�/�/�/�/P/1?�C?�~3}�ɱ ��ߎ?�<��v��?�?��?�~?Oז5AA���SPHERE 2~���/vO�/ �O�O�O�O?�O__ �/<_�O5_r_Y_�_�O �O�_�_%_�_�_�_8o�o\oCo�_�o�oT=ZZ�� �ږ