��  Ij�A��*SYST�EM*��V9.3�0162 9/�2/2021 �A   ����SBR_T �  | 	$SV�MTR_ID � $ROBOT�9$GRP_�NUM<AXIS�Q6K 6NFF~3 _PARAMF�	$�  �,$MD SPD_[LIT  &2*�� � �����$$CLASS ? ���������� VERS�ION�  1r�$' � 1 � T����R-2�000iC/12�5L���  �aiSR22/4�' 80A��
�H1 DSP1-�S1��	P01�.009,  �	�  ���]�   ��# ������������
=��r�9  :!�a������ @H+ � ����?� Y�� �v# < �����  �����&  2��&���>A����$j�?��
"�����&��� )� 	���� ������������� ��A�����y���{����B� U K ���� �5 �:?�����'b�
��E/�/�/�/�/��1�?��3?C?�U?g?��37X���=�����J��4�]��<���\��cx�T�p?�?����0B30/3�L2^2fx��o���������~��%�����8 l�� ^�o�@����� ��*�*�����c	v� 5F���;������Y|��+��\, & ��/�� �8$P�?�������\'%���R��r(��c9	`D� 0��� ����#p�"@��x��Ou_�_�_�_3��_ ?�_��_o��Z���5�Y
��@��p����
��8m� �8u�����pG�Toso�4��?0�?T3^�R"O4OFK��bZOlO~G����H��4�4ٰ�K|4D	 =���,���ܿo(+ ] , " �Bu�O������\'
���h�q��-r(�6_H_Z_#�5�G�Y��-|h��_���� ŏ o�����1��o��o B10J4�Q4^4�o�m:�����(�����2�`8	���� 0��� ������wyF�''nq���`#�5���-�p�/�� l8$�E��s����X��1���E	t����@��5P�!f �<�#S �u��#'  �
�֯�����	01�D;���fF�k� }�������ſ׿�D��V� j�T5^5��������Ɵ؟��x��'��������������+ ��\�O`:"�D�n���[X}�����R
��7e✥�����ʯ�ߥ߷����-
( ��H���#�5�G�Y�k�`}������ "ϊT6^6F�X�j����r�ϔ�����	�������Ϣ����>0 �������
SM #\'	���X��	��r!��h�z��� Ugy�3���� ����"4F�X�������Z��nn���	������/ /&/8/J/\/n/�/�/ �/�/�/�/�/�/?"?2<�2?V?h?z?�?�? �?�?�?�?�?
OC� ~(O����O�O�O �O�O�O�O__0_B_ T_f_x_�_�_�_�_�_ �_@?oo,o>oPobo to�o�o�o�oOJO<O `OrO:L^p� ������ �� $�6�H�Z�l�~����_ ��Ə؏���� �2� D�V�h�z��o���� 0��
��.�@�R� d�v���������Я� ����*�<�N���r� ��������̿޿�� �&�8ϴ���P�ʟܟ ����������"� 4�F�X�j�|ߎߠ߲� ���������h�0�B� T�f�x�������� ��@�r�d�-��Ϛ�b� t��������������� (:L^p� ������  $6HZl~�� ����4�F�X� /2/ D/V/h/z/�/�/�/�/ �/�/�/
??.?@?R? d?v?��?�?�?�?�? �?OO*O<ONO`O� �xO�//�O�O_ _&_8_J_\_n_�_�_ �_�_�_�_�_�_o"o 4o�?Xojo|o�o�o�o �o�o�o�ohO�O�O U�O�O����� ����,�>�P�b� t���������Ώ��<o ��(�:�L�^�p��� ������ʟ&��\ n�H�Z�l�~����� ��Ưد���� �2� D�V�h�z�������¿ Կ���
��.�@�R� d�vψ�������,� >���*�<�N�`�r� �ߖߨߺ�������� �&�8�J�\︿��� ������������"� 4����ϴ�}����ϲ� ��������0B Tfx����� ��d�>Pb t������� N�/
/������p/�/ �/�/�/�/�/�/ ?? $?6?H?Z?l?~?�?�? �?�?"�?�?O O2O DOVOhOzO�O�O�O,/ /�OB/T/f/._@_R_ d_v_�_�_�_�_�_�_ �_oo*o<oNo`oro �o�?�o�o�o�o�o &8J\�O�O�O � __����"� 4�F�X�j�|������� ď֏�����0��o B�f�x���������ҟ �����v?�2�� ��������ί�� ��(�:�L�^�p��� ������ʿܿ�J�� $�6�H�Z�l�~ϐϢ� ������T�F���j�|� ��V�h�zߌߞ߰��� ������
��.�@�R� d�v��������� ����*�<�N�`�r� ��������(�:� &8J\n�� ������" 4FX��j��� ����//0/B/ ��g/Z/�������/�/ �/�/??,?>?P?b? t?�?�?�?�?�?�?�? OOr:OLO^OpO�O �O�O�O�O�O�O _|/ n/_�/�/�/~_�_�_ �_�_�_�_�_o o2o DoVohozo�o�o�o�o �o0O�o
.@R dv���_:_,_ �P_b_*�<�N�`�r� ��������̏ޏ��� �&�8�J�\�n����o ����ȟڟ����"� 4�F�X�j������� � ������0�B� T�f�x���������ҿ �����,�>Ϛ�b� tφϘϪϼ������� ��(ߤ���@ߺ�̯ ޯ�߸������� �� $�6�H�Z�l�~��� ����������X� �2� D�V�h�z��������� ��0�b�T�xߊ�R dv������ �*<N`r �������/ /&/8/J/\/n/�/�/ ���/�/$6H?"? 4?F?X?j?|?�?�?�? �?�?�?�?OO0OBO TOfO��O�O�O�O�O �O�O__,_>_P_�/ �/h_�/�/?�_�_�_ oo(o:oLo^opo�o �o�o�o�o�o�o  $�OHZl~�� �����X_�_|_ E��_�_z������� ԏ���
��.�@�R� d�v���������П, ���*�<�N�`�r� ���������߯үL� ^�p�8�J�\�n����� ����ȿڿ����"� 4�F�X�j�|ώ�ꟲ� ����������0�B� T�f�x���毐�
�� .�����,�>�P�b� t����������� ��(�:�L���p��� ������������  $�߲ߤ�m���ߢ ����� 2 DVhz���� ���T�
/./@/R/ d/v/�/�/�/�/�/�/ >?�/t��`?r? �?�?�?�?�?�?�?O O&O8OJO\OnO�O�O �O�O/�O�O�O_"_ 4_F_X_j_|_�_�_? ?�_2?D?V?o0oBo Tofoxo�o�o�o�o�o �o�o,>Pb t�O������ ��(�:�L��_�_�_ ���_oʏ܏� �� $�6�H�Z�l�~����� ��Ɵ؟���� �| 2�V�h�z�������¯ ԯ���
�f�/�"��� ������������п� ����*�<�N�`�r� �ϖϨϺ�����:�� �&�8�J�\�n߀ߒ� �߶���D�6���Z�l� ~�F�X�j�|���� ����������0�B� T�f�x����������� ����,>Pb t����߽�*�� (:L^p� ������ // $/6/H/��Z/~/�/�/ �/�/�/�/�/? ?2? �W?J?����?�? �?�?�?
OO.O@ORO dOvO�O�O�O�O�O�O �O_b/*_<_N_`_r_ �_�_�_�_�_�_�_l? ^?o�?�?�?no�o�o �o�o�o�o�o�o" 4FXj|��� � _����0�B� T�f�x������_*oo �@oRo�,�>�P�b� t���������Ο��� ��(�:�L�^�p�� ������ʯܯ� �� $�6�H�Z����r�� ���ؿ���� �2� D�V�h�zόϞϰ��� ������
��.ߊ�R� d�v߈ߚ߬߾����� �����0謹�� ο����������� �&�8�J�\�n����� ����������H�" 4FXj|��� � �R�D�h�z�B Tfx����� ��//,/>/P/b/ t/�/�/���/�/�/�/ ??(?:?L?^?p?�? ��?�?&8 OO $O6OHOZOlO~O�O�O �O�O�O�O�O_ _2_ D_V_�/z_�_�_�_�_ �_�_�_
oo.o@o�? �?Xo�?�?�?�o�o�o �o*<N`r �������� �p_8�J�\�n����� ����ȏڏ�Hozolo 5��o�oj�|������� ğ֟�����0�B� T�f�x���������� ү����,�>�P�b� t��������Ͽ¿<� N�`�(�:�L�^�pς� �Ϧϸ������� �� $�6�H�Z�l�~�گ�� ����������� �2� D�V�h��ֿ����� �����
��.�@�R� d�v������������� ��*<��`r ������� p���]���� ������/"/ 4/F/X/j/|/�/�/�/ �/�/�/D�/?0?B? T?f?x?�?�?�?�?�? .�?�?dv�PObO tO�O�O�O�O�O�O�O __(_:_L_^_p_�_ �_�_?�_�_�_ oo $o6oHoZolo~o�oO �?�o"O4OFO 2 DVhz���� ���
��.�@�R� d��_��������Џ� ���*�<��o�o�o ���o�o��̟ޟ�� �&�8�J�\�n����� ����ȯگ����l� "�F�X�j�|������� Ŀֿ���V��ό� ����xϊϜϮ����� ������,�>�P�b� t߆ߘߪ߼���*��� ��(�:�L�^�p�� ����4�&���J�\� n�6�H�Z�l�~����� ���������� 2 DVhz��߰� ���
.@R d��������� �//*/</N/`/r/ �/�/�/�/�/�/�/? ?&?8?�J?n?�?�? �?�?�?�?�?�?O"O ~GO:O����O�O �O�O�O�O__0_B_ T_f_x_�_�_�_�_�_ �_�_R?o,o>oPobo to�o�o�o�o�o�o\O NO�orO�O�O^p� ������ �� $�6�H�Z�l�~����� ��o؏���� �2� D�V�h�z����o ՟0B
��.�@�R� d�v���������Я� ����*�<�N�`��� r�������̿޿�� �&�8�JϦ�o�b�ܟ � ����������"� 4�F�X�j�|ߎߠ߲� ����������z�B� T�f�x�������� �������v� ��Ϭ� �φ������������� (:L^p� �����8�  $6HZl~�� ��B�4��X�j�2/ D/V/h/z/�/�/�/�/ �/�/�/
??.?@?R? d?v?�?��?�?�?�? �?OO*O<ONO`OrO ��O�O//(/�O_ _&_8_J_\_n_�_�_ �_�_�_�_�_�_o"o 4oFo�?jo|o�o�o�o �o�o�o�o0�O �OH�O�O�O��� ����,�>�P�b� t���������Ώ��� �`o(�:�L�^�p��� ������ʟܟ8j\ %���Z�l�~����� ��Ưد���� �2� D�V�h�z�������� ¿���
��.�@�R� d�vψϚ����ϲ�,� >�P��*�<�N�`�r� �ߖߨߺ�������� �&�8�J�\�n�ʿ�� ������������"� 4�F�X�����p����� �������0B Tfx����� ��,��Pb t������� /`�����M/�����/ �/�/�/�/�/�/ ?? $?6?H?Z?l?~?�?�? �?�?�?4�?O O2O DOVOhOzO�O�O�O�O /�O�OT/f/x/@_R_ d_v_�_�_�_�_�_�_ �_oo*o<oNo`oro �o�o�?�o�o�o�o &8J\n��O �O�_$_6_��"� 4�F�X�j�|������� ď֏�����0�B� T��ox���������ҟ �����,���� u�������ί�� ��(�:�L�^�p��� ������ʿܿ� �\� �6�H�Z�l�~ϐϢ� ��������F���|� ����h�zߌߞ߰��� ������
��.�@�R� d�v�������� ����*�<�N�`�r� ������$����:�L� ^�&8J\n�� ������" 4FXj|��� ����//0/B/ T/�������/��
�/ �/�/??,?>?P?b? t?�?�?�?�?�?�?�? OO(O�:O^OpO�O �O�O�O�O�O�O __ n/7_*_�/�/�/�_�_ �_�_�_�_�_o o2o DoVohozo�o�o�o�o �o�oBO
.@R dv�����L_ >_�b_t_�_N�`�r� ��������̏ޏ��� �&�8�J�\�n����� �� ȟڟ����"� 4�F�X�j�|��
�� ů �2�����0�B� T�f�x���������ҿ �����,�>�PϬ� bφϘϪϼ������� ��(�:ߖ�_�R�̯ ޯ�������� �� $�6�H�Z�l�~��� �����������j�2� D�V�h�z��������� ������t�f��ߜ� ��v������ �*<N`r �����(��/ /&/8/J/\/n/�/�/ �/ 2$�/HZ"? 4?F?X?j?|?�?�?�? �?�?�?�?OO0OBO TOfOxO��O�O�O�O �O�O__,_>_P_b_��%�$SBR2 �1�%�P T�0 � �C�/�' �_�_�_�_o o&o8oJo\ono�o�o�o�o�Q�o�_�o '9K]o�� �����o��o#� 5�G�Y�k�}������� ŏ׏�����1�� U�g�y���������ӟ ���	��-�?�"�c� F���������ϯ�� ��)�;�M�_�q�T� ��x���˿ݿ��� %�7�I�[�m�ϑϣ���~i_�������� '�9�K�]�o߁ߓߥ� �����ظ���
��.� @�R�d�v����� ����������*�<�N� `�r������������� ��&
��\n �������� "4FX<f� ������// 0/B/T/f/x/�/n�/ �/�/�/�/??,?>? P?b?t?�?�?�?�?�/ �?�?OO(O:OLO^O pO�O�O�O�O�O�O�O �?_$_6_H_Z_l_~_ �_�_�_�_�_�_�_o  o_DoVohozo�o�o �o�o�o�o�o
. @R6ov���� �����*�<�N� `�r���h����̏ޏ ����&�8�J�\�n� ����������ڟ��� �"�4�F�X�j�|��� ����į֯��̟�� 0�B�T�f�x������� ��ҿ������>� P�b�tφϘϪϼ��� ������(�:��^� p߂ߔߦ߸�������  ��$�6�H�Z�l�P� �������������  �2�D�V�h�z����� ����������
. @Rdv���� ����*<N `r������ �/�&/8/J/\/n/ �/�/�/�/�/�/�/�/ ?"?4?/X?j?|?�? �?�?�?�?�?�?OO 0OBOTO8?J?�O�O�O �O�O�O�O__,_>_ P_b_t_�_jO|O�_�_ �_�_oo(o:oLo^o po�o�o�o�o�_�o�o  $6HZl~ �������o�  �2�D�V�h�z����� ��ԏ���
�� � @�R�d�v��������� П�����*�<�N� 2�r���������̯ޯ ���&�8�J�\�n� ��d�����ȿڿ��� �"�4�F�X�j�|ώ� �ϲϖ��������� 0�B�T�f�xߊߜ߮� ����������,�>� P�b�t������� ���������:�L�^� p���������������  $6�,�l~ �������  2DVhLv� �����
//./ @/R/d/v/�/�/~�/ �/�/�/??*?<?N? `?r?�?�?�?�?�?�/ �?OO&O8OJO\OnO �O�O�O�O�O�O�O�O �?"_4_F_X_j_|_�_ �_�_�_�_�_�_oo 0o_Tofoxo�o�o�o �o�o�o�o,> PbFo����� ����(�:�L�^� p�����x��ʏ܏�  ��$�6�H�Z�l�~� ��������������  �2�D�V�h�z����� ��¯ԯ�ʟܟ�.� @�R�d�v��������� п�������&�N� `�rτϖϨϺ����� ����&�8�J�.�n� �ߒߤ߶��������� �"�4�F�X�j�|�`� ������������� 0�B�T�f�x������� ��������,> Pbt����� ���(:L^ p�������  //�6/H/Z/l/~/ �/�/�/�/�/�/�/?  ?2?D?(/h?z?�?�? �?�?�?�?�?
OO.O @OROdOH?Z?�O�O�O �O�O�O__*_<_N_ `_r_�_�_zO�O�_�_ �_oo&o8oJo\ono �o�o�o�o�o�_�o�o "4FXj|� �������o� 0�B�T�f�x������� ��ҏ�����,�� P�b�t���������Ο �����(�:�L�^� B���������ʯܯ�  ��$�6�H�Z�l�~� ��t���ƿؿ����  �2�D�V�h�zόϞ� ���Ϧ�����
��.� @�R�d�v߈ߚ߬߾� ���������*�<�N� `�r��������� ������
�J�\�n� ���������������� "4F*�<�|� ������ 0BTfx\�� ����//,/>/ P/b/t/�/�/�/��/ �/�/??(?:?L?^? p?�?�?�?�?�?�?�/  OO$O6OHOZOlO~O �O�O�O�O�O�O�O_ �?2_D_V_h_z_�_�_ �_�_�_�_�_
oo.o @o$_dovo�o�o�o�o �o�o�o*<N `rVo����� ���&�8�J�\�n� �������ȏڏ��� �"�4�F�X�j�|��� ����ğ�������� 0�B�T�f�x������� ��ү���ڟ�,�>� P�b�t���������ο ����(��6�^� pςϔϦϸ�������  ��$�6�H�Z�>�~� �ߢߴ����������  �2�D�V�h�z��p� ����������
��.� @�R�d�v��������� ������*<N `r������ ���&8J\n �������� /"/F/X/j/|/�/ �/�/�/�/�/�/?? 0?B?T?8/x?�?�?�? �?�?�?�?OO,O>O PObOtOX?j?�O�O�O �O�O__(_:_L_^_ p_�_�_�_�O�O�_�_  oo$o6oHoZolo~o �o�o�o�o�o�_�o  2DVhz�� �����
��o.� @�R�d�v��������� Џ����*�<�N�