��   v��A��*SYST�EM*��V9.3�0162 9/�2/2021 �A   ����UI_CONF�IG_T  �x L$NUM_�MENUS  y9* NECTCRECOVER>�CCOLOR_C�RR:EXTST�AT��$TOP�>_IDXCME�M_LIMIR$DBGLVL��POPUP_MA�SK�zA  �$DUMMY7]3�ODE�
4CWFOCA �5C+PS)C��g �HAN� � TI�MEOU�PIPESIZE � �MWIN�PAN�EMAP�  ܕ � FAVB ?�� 
$HL�_D�IQ?� qEL3EMZ�UR� l�� Ss�$HMMI�RO+\W �ADONLY� ��TOUCH�P{ROOMMO#{?$�ALAR< ~�FILVEW�	ENB=%%fzC 1"USER:)oFCTN:)WI�u� I* _ED�|l"V!_TITL� �1"COORD�F<#LOCK6%�$F%�!b"EBFOAR�? �"e&
�"�%�!BA�!j ��!�BG�#�!hINS�R$IO}7P}M�X_PKT?$IHELP� {ME�#BLNKC=�ENAB�!? SI?PMANUA�L48"="�BEEY?$X�=&q!EDy#M0qIP0q!�JWD��D7�DSB�� G�TB9I�:J�<ST]Yf2$Iv!_G�v!k FKE�FH�TML�_NAM�#DIMC4:1]ABRIGH83s oD�J7CH92%!FEL0T�_DEVICg1�&USTO_@ � t @ARN$@PIDD�BC�Dn*PAG� ?hA��B�ISCREuE�F���GN�@$�FLAG�@  �&�1  h 	�$PWD_ACC#ES� MA�8��hS:1�%)$LA{BE� $Tz �jHP�3�R�	\} &USRVI >1  < `�Rp*�R��QPRI��m� t1�PTRI�P�"m�$$CL�ASP ����a��R��R `\ S�I�	g ? 1r�$'2 ����R	_ ,��?*���aa1`jbed�`a���� �  ?�C �o��
 �� a�o�o�o%7 �o\n���� E����"�4�� X�j�|�������ďS� �����0�B�яf� x���������O���� ��,�>�P�ߟt��� ������ί]���� (�:�L�ۯp��������ʿܿa`TPTX���l���� s �鶄��$/softpa�rt/genli�nk?help=�/md/tpmenu.dg޿xϊ�ȜϮ�g�&C�U�pwdd�����1�f�U� g�yߋߝ߯�>����� ��	��-����c�u�`��������a��`��b��dc��($R������6�!�Z���ada��c���c��~�N����c����d�a�aJ�  �d]	H�������p���a���`  ���|H Gp��JJ#J�Ffbc :c�B 1)hR �\��_�� �REG VE�D?���who�lemod.ht}m�	singl��doub�tripbrows3b�i {�W������"/����dev�.s�lo/� 1r,	t�/A�//K/ �/�/?�/5?G?Y?k?}?�?� ��?�? �?�?OO+O=OOOaO jE2P�?�O�OqO�O�O �O�E�	�?�?_/_A_ S_e_w_�_�_�_�_�_ �_�_oo+o=oOoao /'yoso�o�o�o�o�o �o1CUgy �������? � 2�D�V�h�z������� �O���Ǐُ.�@� �O	_���������П ˟ݟ���%�7�`� [�m���������oկ ϯ���!�3�E�W�i� {�������ÿտ��� ��/�A��|ώϠ� ������������� B�T�#�5ߊߜ�S�e� K��������,�'�9� K�t�o������� ������߯1�+�Y� k�}������������� ��1CUgy ��k����  2DVhzuߞ� ������ߧ@/ ;/M/_/�/�/�/�/�/ �/�/�/??%?7?`? [?m?;��?�?�?�?�? �?�?O!O3OEOWOiO {O�O�O�O�O�O�O�O �4_F_X_j_|_�_�_ �_�_�_��_o�_�_�BoTobj�$UI_�TOPMENU �1-`�a?R 
d�aQ�)*defau�lt_ ]*level0 *[�	 �o�0�o��o�o	rtpio[�23]�8tpst[1=xY�o��o�=h58e01_l.png�~�6menu5�y�p�q13�z�r�z�t14�{��q��?�f� x���������RT�������1�C�҄p�rim=�qpag�e,1422,1 J���������˟֏�@��%�7�I�ؖ^�class,5R�@��������ϯڔf�13֯��0�B�T�ۓ^�53p�����P��ƿؿۓ^�8� �%�7�I�[�ڟϑ� �ϵ�����Y�`�a �o��mΙq�;�Y��CvtyN}6Hqmf�[0PN�	��c[g164=w��59=x �q)�o���x2��} Q����w�{��O�� ����� ��$�o�H� Z�l�~�����1�����@���� ��e�22 gy���>p�� �	-����n@����e�w�1��@�//*/</��^�?ainedi	�s/��/�/�/�/��co�nfig=sin�gle&^�wintpj��/??*?<? Z�a��J?v?�e~?� �?�?�?�?�?OO 1O�?=OgOzO�O�O�O �O�O�OC�_._@_R_ d_v_�_���_�_�_�_ �_o�_*o<oNo`oro �oo�o�o�o�o�o �o8J\n�� !������� "�F�X�j�|�����/� ď֏�������B�@T�f�x������N�� ҟ�/�UE��O���As��:�_���G�u�� ���n�l�2��V��h�L�:�6G�u7� �����ÿտ�2� ��/�A�S�e����π�ϭϿ��������"�1�/�A�S�e�w� �ϛ߭߿������߄� �+�=�O�a�s��� �������������6
�?�Q�c�u����$��74�����������V<��>�5	TP?TX[209��^DY24��,��d�Y18~���at0�2��aA��=��tvB�4FX.�0p-1pi�S:��$treevie�w�#��3��&du�al=o�81,26,4�1/C/U/ �y/�/�/�/�/�/b/��/	??-???Q?��;���53/$���? �?�?�/OO)O;OMO _O�?�O�O�O�O�O�OHd?v?��1�?$2��8H_Z_l_ �6�O��edit�� _2_�_ �_�_������_�S�_ Qocouo$vo�o핪o #�o��o�o1 CUz�os��� ���
��y�3�Z� l�~�������sO؏� ��� �2���V�h�z� ������?����
� �.�@�ϟd�v����� ����M������*� <�˯N�r��������� ̿[����&�8�J� ٿnπϒϤ϶���wo �o�ϭo"߉'�E�W� i�{ߎߟ߱���1��� ����/�A�S�e�w� 9������������� e�>�P�b�t�����'� ����������: L^p���5� �� $�HZ l~��1��� �/ /2/�V/h/z/ �/�/�/?/�/�/�/
? ?.?����d?߈?�� ��?�?�?�?�?OO )O�?5O_OqO�O�O�O �O�O�O��_&_8_J_ \_n_�_�/�_�_�_�_ �_�_�_"o4oFoXojo |oo�o�o�o�o�o�o �o0BTfx� ������� ,�>�P�b�t�����'� ��Ώ�������:� L�^�p�����C?U?ʟ y?�UO�O�#�5�G� Y�k�~�������ůׯ �����1�C�_z� ������¿Կ��
� �.�@�R�d��Ϛ� �Ͼ�����q���*� <�N�`���rߖߨߺ� ��������&�8�J� \�n��ߒ������� ��{���"�4�F�X�j� |�������������������*defa�ult؞*level8a���Y��w�! tp�st[1]�	�y��tpio[23���u�d��,>menu7�_l.pngA&^13cp5x]4�[4�u6cp� ��	//-/?/��c/ u/�/�/�/�/L/�/�/�??)?;?M?�"p�rim=^pag?e,74,1R?�?��?�?�?�?�"f6class,13�?�OO0OBOTO�?�25�ZO�O�O�O�O�O�# �<~O_$_6_H_Z_]?o218v?�_�_�_�_�_�O�26�_o-o?o�QocoB�$UI_�USERVIEW� 1�����R 
�� jo䒞o�o=m�o�o 	-?�ocu� ��N����� �o$�6�H�������� ��ˏn����%�7� I��m��������`� ԟ�X�!�3�E�W� i��������ïկx������/�A��*�zoomT�ZOOMIN�S�񯺿 ̿޿�ϥ�&�8�J� \�n�ϒϤ϶������<*maxres~n�MAXRES�� �ω�R�d�v߈ߚ�=� ����������*�<� N�`�r�߃���� ������&�8���\� n�������G������� ����3A��| ����g�� 0B�fx�� �Y���Q/,/ >/P/b//�/�/�/�/ �/q/�/??(?:?� K?Y?k?�/�?�?�?�? �? O�?$O6OHOZOlO O�O�O�O�O�O�?�O �O	_{OD_V_h_z_�_ /_�_�_�_�_�_
o�_ .o@oRodovoa