��   !��A��*SYST�EM*��V9.3�0162 9/�2/2021 �A   ����BIN_CFG�_T   X �	$ENTRIE�S  $Q0�FP?NG1F1*O2F2OPz ?�CNETG  ��DHCP_CTR�L.  0 �7 ABLE? $�IPUS�RET�RAT�$SE�THOST��N�SS* 8�D��FACE_NU�M? $DBG_�LEVEL�OM�_NAM� ! ���* D �$PRIMAR�_IG !$AL�TERN1�<W?AIT_TIA �� FT� =@� LOG_8	��CMO>$DN�LD_FI:�S�UBDIRCAP� ��8 .� 4� H�A�DDRTYP�H NGTH��Y�z +LS�&$ROBOT2�PEER2� MA�SK4MRU~O�MGDEV�$D�PINFO�m $$$X�A�RCM�T A$| ��Q�SIZ�X�� T�ATUSWMAI�LSERV $�PLAN� <$�LIN<$CLyU���<$TO�oP$CC�&FR�&��JEC�!�%E�NB � ALA5R�!B�TP�/3�V8 S��$VkAR79M ON,6���,6APPL,6P�A� -5B +7POR���#_12ALE�RT�&�2URL �}�3ATTA�C��0ERR_T7HRO�3US�9�!��8R0CH- YDM�AXNS_�1��1AMOD�2AI�� o 2A� (1APoWD  � LA ��0�ND)ATRYsFDELA�C2@�'`AERSI�1A�'�RO�ICLK�HM8t0�'� XML+ \3_SGFRM�3T� fXOU�3Z G_��COPc1V�3Q�'qC�2-5R_AU�� � XRN1oUPD�XPCOU�!SF�O 2 
$�V~Wo�@YACCܳH�QSNAE$UM�MY1�W2?N��RDM*	� $�DISc �SM}B�
 T �	BCl@DCI2�AI&P6EXPS��!�PAR� `R{ANe@  ��QCL� <�(C�0�SPTM
U� PWR�-hCf��SMo l5��!�"%�7Y�P"�% 0�fR�0�e=P� _DLV�De&�SNo3 
j��hX_!`�#Z_I�NDE,C_pOFF,� ~URnyD�  �*s�   ts �!pMON�r�sD��rHOU�#�EyA�v�q�v�q�vL�OCA� Y$Nާ0H_HE��rPI"/  d	`GARP�&�1F�#W_~ �I!Fap;�FA�D�01#�HO�_� �R�2P$`�S�wTEL	% P dK  !�0WO�`� �QE� LV��k�2H#ICEدڀ�P�$d�  ��������
���
��`S$Q���  1rc�$'0 �
����F����"�S�L���$� 24� ������e��� 4����! �ʟ����-�4�Ɵ��8�I�L����p_V`4�� S�z�������¯ԯ毀��
��.�@��� _?FLTR  �?�W �������!�ޛnx4�2ޛ8�{SHE`D 14�E P'��I�ٿ ��:���^�!ς�E� ��iϷ��ϟ� ���$� ��H��l�/�Aߢ�e� �߉��߭������D� �h�+��O��s�� ����
���.���R�� ^�9�����o������� ����<��r5 �Y�}��� �8�\�Cy�������PP�P_L�A1e�x/!1.9"0/��8%1I/�2551.�%@/��Q�7#2>/P.� d/v/�/�/�&3�/P.-0�/�/ ??�&4.?P.�0T?f?x?�?�&5�?P.@�?�?�?O�&6OP.�@�DOVOhOzOT�aP����(���Ӱ��� OQ� ��N<0_ e_w_J_�_�_�_�_�_�_�P�_%o7oIoo moo�o�obo�o�o�o��N�o�T�5 |�
ZDT Status�oD�����}iRCon�nect: ir�c�t//alertb~���+��wt�Y�k�}��������2A�P�RJ������  ��$�6�H�Z�l�~��������ƟQs$$c�962b37a-�1ac0-eb2�a-f1c7-8�c6eb579e?ef5  (H��@l=�O�a�s���A
��X�'R��)z��� *t��2u+Q!T,$4�񯨰*!߯�� @�'�M�v�]������� п����ۿ����N��5�r�Y������&%PDM_Q	�&+"SMB 
 &%U�#l��O����� Iߌ�� �'��_CLN�T 2&)9�4+t	�|�#|j߯ߎ� ������������Q� 0�u��f�������
.SMTP_CT�RL R� P% ��4�	t��"�c���R� ��v���#|��N�Q��΢��7������ S��US?TOM ����&P �TT�CPIP�����'xU"Ri EL$�&%#Q� H!T�т��rj3/_tpd�� + ��?!KCL��������!CRT�.uR�!OCONSv�
�ib_smon~r