��   #��A��*SYST�EM*��V9.3�0162 9/�2/2021 ?A   ������DMR_SH�FERR_T �  $OF�FSET  � 	j/GRP�: $M�A��R_DONE�  $OT_�MINUSJ  �	sPLzdCO{UNJ$REFj�PO{��I�$BCKLSH_�SIG�EAC�HMSTj�SP9C�
�MOVn ~�ADAPT_IN�ERJ FRI}CCOL_P,=MGRAV��� HISIDS�Pk�HIFT_Z7 O �Nm��MCH� S�ARM_PARAOw dcANGo �y2�CLDE|7�CALIB�Dn$GEARr�2(�� �RING��<$r]_d�REL3�� 1  	K�\�CLo:o � �AX{ � $PS_�T�I���TIME� �J� _CMYD��"FB�VS >�&CL_OV�� oFRMZ�$DE�DX�$NA� =%�CURL�qW���TCK5��FMSV>�M_LIF	���;8G:w$�A9_0M:_��=�93x6W�� �"�PCCOM,��FB� M�0�oMAL_�ECI��PL!�"DTY�kR_�"�5L#�1E�NDD��o1� �5M�  ��PL� W ��  $STAL#T�RQ_M��0K$N}FS� �HY�J� *|GI�JI�JI�E#�3AnCuB�A�E��$�ASS> �S��	Q�����@�VERSI� W�  1r��$S 1'X_ ���M@���n_Y_�_}U����N@�1T���<���h� ƅ7��X_�_�_ �_x]2P+b3oz[QTo�Bl��J�Ο�s 21��?�����k;Ao�o=ogl�o�o�o�t� 7u�gB@Mv Ww#�o�s���d���<���=L���.�3?�/���@�O�t� ��������Ώ����0�(�:�� 	Ue�ps�]���T  2� ğ֟�����0�B�T�f��R�������� Ưد���� �2�D� V�h�z�������¿Կ ���
��.�@�R�d� vψϚϬϾ������� ��*�<�N�`�r߄� �ߨߺ��������� &�8�J�\�n������<��������� &�8�J�\�n������|(���������� 2/hS�w�`����
�$&4� 1D\��O�Z�HJUI�¡�M$x�L?�Y�L!GP��L��$O�:��OU��I�٭�J�NI�x��B�  ��B���@o����@B�bD��g��ӽk��H�)N�>�N���Hx���I��G�ɽ�~8�/�>�JI¦�J��N�R�U�VoJO�g/��/v/�/�T��U��}T�!�$^�^�^��^���U� �� CPV;^��B$��BI�h�F�yB�cc�,������+~$���02�Fx/�0��,�&0���-<�ɾ�`��A[�>���d�3���Q��^ �]�%�APPRO�0PAcRT�/V�� ���S�2,3yBI���G�B�a��,�}����>*?s1BIܲ��G6�0y�,������BR>��]����A�Z:>�Ε�/��%:w?�?�?�? ����8:3h{B�I��G�]B��[@�,�/����z�?h��@O��G�C�@�@����d�/  ���`pA6�>�Ɩ��8�K��&��:OLO^O�=�uF\� 0AN5Ir���"���n��:�B�`Y�?��C'`b�OR��j��R��;�h�B�Wx��nC'L��M>�/Y�q�A��r4?J{q��S�?�-R�_A  �RP�_PALLOAD<+_U�  ��!EU��C�������:�SB�h������C'b��j_�������;s�^P�����fC'S��M;������lVA��
�?Y9-�&?K.>ߞ��_�_��_T�)0�4BWP;�NS�t��s$��9�r`A���?C'm`*o�������9�h�`/��RC'�i�R>nsz����ZA�χ?.��e�*9�=ċC�R�U�o�oR��|�Ip�DAU�3��BJV�E��iB�T��,��{��SɪO�_�BJ�E����p&�,���p��R>%߾�`\�A��>����6/�O�!__��<��x�3��BJ�F��B�S �@����Z�c/:��V����F ^�w�,��f�)n;æ������A9�~.CHS;���

��.��;�x��3v�BJ���F�[B�Q1�,����d�j��m`BJ'�F��`B�R�,��y��f�R>���O�� A�->Çb�.��;�ʏ܏�^BVB}o�%���BJ����p�B�+�+�Iy�K�I~%���֐���&e�B� ��*�k��6�:R> e�������:,�A�J���v��1i���P��&TtUN[��$��GQ�O��NS^_����Y�ʃB������.C)�}J�oU���������B���%����C)D�ޒ^��{�;��A���@���Y��@�Ma<��K_��m,9�����NSt���M�����B�l}
p�C)���pm��R���	B�[����C)�G�^a�ue�}A�� 9?���?��@tb�����0�-,��0n���!A��CA�ҧ���K0B��u�5g��חf�M��A��wx���OB��|4"�T��r���M:C����I��Al�?N��r��0��:�̶TTAUGHTPOU������=��IA�S���W�B�z��4Y��V��*��oA�M!��OnB�}"��~���~����'��A\��?I?�*���^8O���Ϯϳ��������π�"�4�F�X�)���0oJ��B����@0���k�B�xd��D'���Л��@��@��[dB��t���K����ԩ�ݾM�C�����Ant)�?Ey̽�	
�=�k�C�� %	>��FAULT�.� 1�B�B�B@��%��ԵB��i��Z3����Q>�k@��A�������?�[��Ɖ`����§�Am"��?(i#��_9�7O������ 1��B�U"��@�����?��-�����!��@�����>����՟h<�ӻ��_����Am$?(E���}�Y���ߌ�ђ�c��2��1Z%����4�B49���._�B�	AS�C��� �B44{�.�K?B��AS�,�C�% � ��y�A+4��>{o>��_ý�^}�����_ASSEMBL�Yk��� A��C �3�;BI�K�E�NB�Y
@�N��*���BI����F	?B��dK�,�k������=�����kA�K>�����Q>���z������>ʎ�&
�
/ ����$PLCL_GR�P 1���;!�� p�R��?�  T+��?y�cT)�/�/ �I�/�/�/�/�/?�/�%??I?4?m??N,z���T"t�?~�=l)