��   
��A��*SYST�EM*��V9.3�0162 9/�2/2021 �A   ����CCLINKR�D_T  4� 9$ASGUO�P  $HD�SHKENB?E�RROR_1PO�ST?WARNI�NGISEQST�=pCPU?IN�_CLR_BIT�S�	WORD?U�SETIMOVR�LM?SCAN_�MODE  ��� �BAUDR�ATE? $� U�LE_ID� $�NUM_STAT�ION? $�_�NO�MAKER�_C� DEVI�CESW_VE;RS�DLE. �� �O5LI�?$REMRE� I�$AO_CH_�� kIrREG_�OUT�_HEA@��� �� �H� O_A_M��B��MIN� <^CV�WAIT�PS_�DAT_���!�TY>_SER�VE_�*$11*L�?!&'L2O+3O+4<�5$I �MvEV�*HBޯTVAL�WD1G���CME�%�$N#�$]#DIAG�N#�!�'l#�!{#�!5z�&6�AUTO
!CHG? �a~<2DUMMY5!1�O5+1  D&C�F/ 4 $�� P_SWITCH�#EBU;1�4�$��1]"��&�! �l>0LOC0NABL��2��Q?1_MASK<2�4SPTJ4Q2�<2�<3�<3�7��8CC:J8HaC�7XTR��6��B�6�1INDEX��#LOCK A ' �6�@�5] �Gl �B�U>!�H�EPROC��A�A�Fp�AZ�A�@��$�@�ASS  �S��<Q��7��71P�5:W  �1r�$' 2� <U7�  ���eP�_�X����U�R #r? 	�V�S
 �P��CQ�W���V720P22 070315�_2��o2o  BR�_ �_Xe a�_�_�_�_opo�o:lkWCFGx0�ZX�P��kWDG 2Mx\��o�T�Rt�����o�� ���xq*�<��`� r���S�����̏ޏe ��&��7�I�[�m� �����ȟ������ ߟ4�F�X�3zv�2�b!u