��   D�A��*SYST�EM*��V9.3�0162 9/�2/2021 �A 
  ����CELLSET�_T   �w$GI_STY�SEL_P }7T  7ISO:iRibDiTRA�R�>�I_INI; �����bU9AR�TaRSRPNS�1Q234�5678�Q
TROBQACKSNO� �)�7�E�S �a�o�zU2 3 4 5 6 7 8awn&GINm'D�&��) %��)4%��)P%�̖)l%SN�{(OU���!7� OPTNAA�73�73.:B<;�}a6.:C<;CK;C�aI_DECSN�A�3R�3�TRY�1��4��4�PTHCN�8D�D�INCYC@HG��KD�TASKOK �{D�{D�7:�E� U:�Ch6�E�J�6�C�6U�J�6O�;0U��:IATL0RHaRbHaRBGSOLA�6�VbG�S�MAx��V�8�Tb@SEGq�Tp��T�@REQ� d�drG�:Mf�GJO_HFAUL�Xpd�dvgALE�  �g�c�g�cvgE� �H<�dvgNDBR�H�dgRGAB�Xtb~���CLMLIy@�   $�TYPESIND�EXS�$$CL�ASS  �S��lq����apVERSIONix�  1Gr�$'61�r���p��q�t+ U�P0 �xS�tyle Select 	  ����r�uReq. /�Echo���yA�ck���sInitiat�p�r�sE�t@�O�a�p����	��  ��*��������:q��������q��sO�ption biGt A��p�B�����C�Decis��cod;��zTr?yout mL���Path seg�J�ntin.�I�I�yc:��Tas�k OK��!�Ma�nual optK.r�pAԖBޟ�ԖC�� decs�n ِ�Robo�t interl�o�"�>� iso)l3��C��i/�"�z�ment��z��ِ����_�stat�us�	MH F�ault:��ߧAler��%��p@r7 1�z L���[�m�+�; LE_COMNT ?�y�   ��䆳� Ŀֿ�����0�B� T�g�xϊϜϮ����� ������,�>�P�b� t߆ߘߪ߼������������U��9r���   ��ENAB  ���u����������ꐵME�NU>�y��NAM�E ?%��(%$*4���D��p2�k�V� ��z����������� ��1U@Rdv ������� *<u`��� �����/;/&/ _/J/f/n/�/�/�/�/ �/?�/%??"?4?F? X?j?�?�?�?�?�?�? �?�=