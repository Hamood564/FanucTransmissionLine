��   ��A��*SYST�EM*��V9.3�0162 9/�2/2021 �A 	  ����DRYRUN_�T  4 �$'ENB  �$NUM_POkRTA ESU@�$STATE }P TCOL_���PMPMCmGR�P_MASKZE�� OTIONNLOG_INFON�iAVcFLTR�_EMPTYd ?$PROD__ L ��ESTOP_D�SBLAPOW_�RECOVAOP�R�SAW_� G� %$INI�T	RESUME�_TYPENDIST_DIFFA $ORN41� 8d =R  �&J�_  4 u$(F3IDX��_ICI  �MIX_BG-yy
_NAMc �MODc_US�d�IFY_TI�� �MKR�-  $L{INc   "o_SIZc_l��� �. h $USE_FL�C 3!�:&iF*SIAMA7#QC#QBn'oSCAN�AX�+�IN�*I��_COUNrRO( ��!_TMR_VA�g#h>�i a �'` ����1n�+WAR�$�iH�!�#N3CH��PE�$O�!PR"�'Ioq7iOq���OoATH-� P $ENA#BL+�0B�T���$$CLA�SS  ����A��5��5�0V�ERS�G  1r�6|/ E5���E����-@]F@AbE��%A�O���O��O����3EI2>K�2_ _2_D_V_ h_z_�_�_�_�_�_�_��_
oo.o�ONV?y"HI@ ���lj�{o�����lj���� � �2>I  4%	IO2CC �K:o�� qT�T�%
CUBE�4���	Csשd%�
SPACECH�EC�o)VUl#j%S�1woAt �������� I�(�:��c$"+ �ktK�-@����bA��X��@A-@vNڏ� ���"�4�F�X�j�|� ��������bFoAǁoA ���
��.�@�R�d� v���������ЯDZM�_��>�C� 2�lǏ1�C�U�g� y���������ӿ��� 	�Ɯ#�<�N�`�rτ� �ϨϺ��������� �8�J�\�n߀ߒߤ� �����������"�-� F�X�j�|������ ��������)�;�T� f�x������������� ��,7�Pbt ������� (:E^p�� ����� //$/ 6/ASl/~/�/�/�/ �/�/�/�/? ?2?D? Ch�4�0��{?��