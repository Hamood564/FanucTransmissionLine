��   ?3�A��*SYST�EM*��V9.3�0162 9/�2/2021 �A   ����MN_MCR_�TABLE  � � $MAC�RO_NAME �%$PROG�@EPT_IND�EX  $O�PEN_IDaA�SSIGN_TY�PD  qk$�MON_NO}PREV_SUBy �a $USER_�WORK���_L� MS�*RTN�   &SO�P_T  �� $�EMGO���RESET��MOT|�HOALl�� 2��STAR PDIU8G9GAGBG�C�TPDS�R�EL�&U� 9�� �EST����SFSP�C����C�C�N	B��S)*$8*$U3%)4%)5%)6%)�7%)S�PNST�Rz�"D�  �$�$CLr   �����!������ VERSION��(  �1r�:LDUI_MT  ��� �����$MAXDSRI� ��5
�$�.1 �%� � d%T{1 f L 1�����%A_TOOcL_P2�?��G����!���!K2SHU�TT?f?x1�2�?�6H*�6�82O52�?�8�Bv?OO 0�4@J�4O1O�?�<J�6��1�3  lose� hand�O�8	 �O_ �"�4-U�@elax�O�OU_{_�*_�Cglogic }_Z_�_~_�]
@�_o �_<o�_�_ro!o�o�o Wo�o�o�o�o�o8 �o5n/�S� w����4��� j����=�O���֏�� ������0�ߏT��� O���K���o������� �,�۟�b����5� G���k���򯡯��(� ׯL����������� g�y�����ӿ� Z�E�~�-�?ϴ�c��� �ϙ��� ���D���� z�)ߞ߰�_ߙ��ߕ� 
����@���=�v�%� 7��[������� �<�����r�!���E� W�����������8 ��\W�S� w���"4� j�=O�s� ���0/�T/// �/�/�/�/o/�/�/�/ ?�/�/?b?M?�?5? G?�?k?�?�?�?�?(O �?LO�?O�O1O�O�O gO�O�O�O_�O�OH_ �OE_~_-_?_�_c_�_ �_�_o ooDo�_o zo)o�oMo_o�o�o�o 
�o�o@�od% _�[���� *�<��%�r�!���E� W�̏{�ɏ���Ï8� �\���������ȟ w�������"�џ�� j�U���=�O�įs�� �����0�߯T��� ��9�����o������� �ɿۿP���Mφ�5� Gϼ�k��Ϗϡ��(� �L���߂�1ߦ�U� gߡ����������H� ��l��-�g��c��� ������2�D���-� z�)���M�_������� 
����@��d% ������ *��%r]�E W�{����8/ �\///�/A/�/�/ w/�/�/�/"?�/�/X? ?U?�?=?O?�?s?�? �?�?O0OOTOOO �O9O�O]OoO�O�O�O _�O�OP_�Ot_#_5_ o_�_k_�_�_�_o�_ :oLo�_5o�o1o�oUo go�o�o�o�o�oH �ol-���� ����2���-� z�e���M�_�ԏ���� �����@��d��%� ��I���П������ *�ٟ�`��]���E� W�̯{�𯟯��&�8� #�\�����A���e� w������"�ѿ�X� �|�+�=�w���s��� �ϩ����B�T��=��
Send Ev�entU�5�SE?NDEVNT��3�{)i� %	}��Data�ߘ�DA�TA�߿���%~}�SysVar�SYSVY��+>1�%Get��Z�OGET��,���%Reques?t Menu����REQMENU!���-��?߀�;ߤ�_� �����������F ��j+�O�� ���0��f xc�K]��� ���>/)/b//#/ �/G/�/k/}/�/?�/ (?�/�/^??�?�?C? }?�?y?�?�?�?$O�? !OZO	OO�O?O�OcO uO�O�O�O _�O�OV_ _z_)_;_u_�_�_�_ �_�_o�_@o�_o;o �o7o�o[omo�o�o �oN�or!3 �W������ 8���n���k���S� e�ڏ����������F� 1�j��+���O�ğs� �������0�ߟ�f� �����K���ү���� ����,�ۯ)�b��#� ��G���k�}���� (�׿�^�ς�1�C� }��ϵ��ϝϯ�$��� H���	�Cߐ�?ߴ�c��u��$MACRO�_MAX:����_��Ж���SOPENBL ?���������r�r�A���PD�IMSK�����Y�SUc�u�TP�DSBEX  -�q�U����n� ���