��   -�A��*SYST�EM*��V9.3�0162 9/�2/2021 �A   ����CELL_GR�P_T   �� $'FRAM�E $MOUNT_LOCC�CF_METHO�D  $CP�Y_SRC_ID�X_PLATFR�M_OFSCtD�IM_ $BAS=E{ FSETC���AUX_ORD�ER   ��XYZ_MAP� �� �L�ENGTH�TTCH_GP_M~ �a AUTORAI�L_4�$$C�LASS  ������D��D�VERSION�  �1r�8LOOR� G��DD<Z$?���q��Mn,  1 <DYX< [�����D'�i�����iO/a/s/A/p�/�/�/$ �/��/�/	;�$MNU�>A>"�  	� <iU{��H[;�u��IW�Ux�< ���d���4'��gEB�Cr�8�SC���?��0=8I0Z�;�t�Q0VU0��< �\0�1a0�je4sm4;u;zQ0��;���J�ӿUw�<��v�f����e0kE���;<C��� ��4i�V�k��K������J�?V�;�;'^}����;������N����)K/C�����i# 5O�-O!/}OcO�O�O �O�O�O�O�O_1_�~5NUM  ��9	a� �0�TOOL%?\ =
;7�;�.AE�Yٿ�T�QÌ��C�[�Y3��.�Q'W����U3�PC�_ 0OBO4Zeo?_goMo oo�o�o�o�o�o�o�o #Q7i�m���SX�QcS[
nY��D