��   (�A��*SYST�EM*��V9.3�0162 9/�2/2021 �A 	  ����PASSNAM�E_T   0� $+ �$'WORD  �? LEVEL � $TI- OU�TT  &F/�� $SET�UPJPROGR�AMJINSTA�LLJY  ?$CURR_O��USER�NUM��STSTOP_TPCHG V oLOG_P NT��N�  6 CO�UNT_DOWN��$ENB_P�CMPWD� $kDV_� IN� �$C� CRE���A RM9� T9DIAG9(�>LVCHK FULLM/�Y{XT�CNTDޏMENU�AU�TO+�FG_D�SP�RLS�U��BURYBAN���GI�VfE�NC/  ~CRYPTE�    ��$$CL( L ����[!�� d P V�� IONX(�K 1r�$DC�S_COD?�|��_%�  W�'q_� �/�(S  Z*%�� \ �&�A9�1�"[!	 
 $b!��= ?4?B?X?f?|?�?�? �?�?�?�?�?OO0Op>OTO���#SUP� � :�VOhO�#F��O�O�O�� C \Q��_ 0��� V�[t�&��j���D �Op_��.W,_��K �V��U�YqILUGH �1[) K �)�_oo/oAo Soeowo�o�o�o�o�o �'�_�o#5GY k}������o ���1�C�U�g�y� ��������ӏ��	� �-�?�Q�c�u����� ����ϟ�����)� ;�M�_�q��������� ˯ݯ���%�7�I� [�m��������ǿٿ ����!�3�E�W�i� {ύϟϱ��������� ��/�A�S�e�w߉� �߭߿��������� +�=�O�a�s���� �������� ��'�9� K�]�o����������� �������#5GY k}������ ��%