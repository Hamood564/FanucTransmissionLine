��   �A��*SYST�EM*��V9.3�0162 9/�2/2021 �A   ����FSAC_LS�T_T   8� $CLNT_�NAME !�$IP_ADDR�ESSB $AC�CN _LVL � $APPP  _V �$8 AO ? ���z�����o VERS�IONw  1r�$'�DEF\ w { �� ���ENA'BLEw �������LIST 1 ��  @!ȁ������ 
[.@�d�� ���/�3//W/ */</�/`/�/�/�/�/ �/�/�/??S?&?8? J?�?n?�?�?�?�?�? O�?�?OO"OsOFO�O jO|O�O�O�O�O_�O �O6__\_B_�_f_x_ �_�_�_�W